
module mul32_3_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n321, n324, n327, n330, n333, n336, n339, n342, n345, n348, n351,
         n354, n357, n360, n363, n366, n369, n372, n375, n387, n390, n393,
         n396, n399, n402, n405, n408, n416, n419, n422, n425, n428, n431,
         n434, n437, n440, n443, n446, n449, n458, n461, n465, n469, n471,
         n473, n475, n477, n479, n481, n483, n485, n487, n489, n491, n493,
         n495, n497, n499, n501, n503, n505, n507, n509, n511, n513, n515,
         n517, n519, n521, n523, n525, n527, n529, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n600, n601,
         n602, n603, n604, n605, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n620, n621, n622, n623, n624, n625,
         n627, n630, n631, n632, n633, n634, n635, n636, n637, n638, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n667, n668, n669, n670, n671, n672, n673, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n714, n715, n716, n717, n718, n719, n721, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n734, n735, n736, n737,
         n738, n739, n744, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n833,
         n835, n836, n838, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n999, n1000, n1002, n1003, n1004, n1005, n1009,
         n1010, n1011, n1012, n1018, n1019, n1020, n1022, n1026, n1028, n1029,
         n1036, n1038, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818;
  assign n321 = a[1];
  assign n324 = a[3];
  assign n327 = a[5];
  assign n330 = a[7];
  assign n333 = a[9];
  assign n336 = a[11];
  assign n339 = a[13];
  assign n342 = a[15];
  assign n345 = a[17];
  assign n348 = a[19];
  assign n351 = a[21];
  assign n354 = a[23];
  assign n357 = a[25];
  assign n360 = a[27];
  assign n363 = a[29];
  assign n366 = a[31];
  assign n465 = b[0];
  assign n469 = b[1];
  assign n471 = b[2];
  assign n473 = b[3];
  assign n475 = b[4];
  assign n477 = b[5];
  assign n479 = b[6];
  assign n481 = b[7];
  assign n483 = b[8];
  assign n485 = b[9];
  assign n487 = b[10];
  assign n489 = b[11];
  assign n491 = b[12];
  assign n493 = b[13];
  assign n495 = b[14];
  assign n497 = b[15];
  assign n499 = b[16];
  assign n501 = b[17];
  assign n503 = b[18];
  assign n505 = b[19];
  assign n507 = b[20];
  assign n509 = b[21];
  assign n511 = b[22];
  assign n513 = b[23];
  assign n515 = b[24];
  assign n517 = b[25];
  assign n519 = b[26];
  assign n521 = b[27];
  assign n523 = b[28];
  assign n525 = b[29];
  assign n527 = b[30];
  assign n529 = b[31];

  XOR2_X2 U319 ( .A(n1042), .B(n1041), .Z(n532) );
  NAND2_X4 U322 ( .A1(n979), .A2(n597), .ZN(n533) );
  NOR2_X4 U324 ( .A1(n1043), .A2(n1046), .ZN(n596) );
  NAND2_X4 U325 ( .A1(n1043), .A2(n1046), .ZN(n597) );
  NAND2_X4 U330 ( .A1(n980), .A2(n602), .ZN(n534) );
  NOR2_X4 U332 ( .A1(n1050), .A2(n1047), .ZN(n601) );
  NAND2_X4 U333 ( .A1(n1050), .A2(n1047), .ZN(n602) );
  XOR2_X2 U334 ( .A(n610), .B(n535), .Z(product[60]) );
  NAND2_X4 U340 ( .A1(n981), .A2(n609), .ZN(n535) );
  NOR2_X4 U342 ( .A1(n1051), .A2(n1056), .ZN(n608) );
  NAND2_X4 U343 ( .A1(n1051), .A2(n1056), .ZN(n609) );
  XNOR2_X2 U344 ( .A(n623), .B(n536), .ZN(product[59]) );
  NOR2_X4 U350 ( .A1(n633), .A2(n617), .ZN(n615) );
  NAND2_X4 U352 ( .A1(n983), .A2(n982), .ZN(n617) );
  AOI21_X4 U353 ( .B1(n982), .B2(n627), .A(n620), .ZN(n618) );
  NAND2_X4 U356 ( .A1(n982), .A2(n622), .ZN(n536) );
  NOR2_X4 U358 ( .A1(n1057), .A2(n1062), .ZN(n621) );
  NAND2_X4 U359 ( .A1(n1057), .A2(n1062), .ZN(n622) );
  NAND2_X4 U366 ( .A1(n983), .A2(n625), .ZN(n537) );
  NOR2_X4 U368 ( .A1(n1063), .A2(n1070), .ZN(n624) );
  NAND2_X4 U369 ( .A1(n1063), .A2(n1070), .ZN(n625) );
  NAND2_X4 U374 ( .A1(n673), .A2(n635), .ZN(n633) );
  NOR2_X4 U376 ( .A1(n656), .A2(n637), .ZN(n635) );
  NAND2_X4 U378 ( .A1(n646), .A2(n984), .ZN(n637) );
  AOI21_X4 U379 ( .B1(n647), .B2(n984), .A(n640), .ZN(n638) );
  NAND2_X4 U382 ( .A1(n984), .A2(n642), .ZN(n538) );
  NOR2_X4 U384 ( .A1(n1071), .A2(n1078), .ZN(n641) );
  NAND2_X4 U385 ( .A1(n1071), .A2(n1078), .ZN(n642) );
  NOR2_X4 U390 ( .A1(n651), .A2(n648), .ZN(n646) );
  OAI21_X4 U391 ( .B1(n648), .B2(n652), .A(n649), .ZN(n647) );
  NAND2_X4 U392 ( .A1(n985), .A2(n649), .ZN(n539) );
  NOR2_X4 U394 ( .A1(n1079), .A2(n1088), .ZN(n648) );
  NAND2_X4 U395 ( .A1(n1079), .A2(n1088), .ZN(n649) );
  NAND2_X4 U398 ( .A1(n986), .A2(n652), .ZN(n540) );
  NOR2_X4 U400 ( .A1(n1089), .A2(n1098), .ZN(n651) );
  NAND2_X4 U401 ( .A1(n1089), .A2(n1098), .ZN(n652) );
  NAND2_X4 U410 ( .A1(n987), .A2(n661), .ZN(n541) );
  NOR2_X4 U412 ( .A1(n1099), .A2(n1110), .ZN(n660) );
  NAND2_X4 U413 ( .A1(n1099), .A2(n1110), .ZN(n661) );
  NAND2_X4 U416 ( .A1(n988), .A2(n664), .ZN(n542) );
  NAND2_X4 U419 ( .A1(n1111), .A2(n1122), .ZN(n664) );
  NAND2_X4 U424 ( .A1(n989), .A2(n669), .ZN(n543) );
  XNOR2_X2 U428 ( .A(n679), .B(n544), .ZN(product[51]) );
  NOR2_X4 U434 ( .A1(n680), .A2(n677), .ZN(n673) );
  NAND2_X4 U436 ( .A1(n990), .A2(n678), .ZN(n544) );
  NOR2_X4 U438 ( .A1(n1137), .A2(n1150), .ZN(n677) );
  NAND2_X4 U439 ( .A1(n1137), .A2(n1150), .ZN(n678) );
  NAND2_X4 U442 ( .A1(n991), .A2(n681), .ZN(n545) );
  NOR2_X4 U444 ( .A1(n1151), .A2(n1166), .ZN(n680) );
  NAND2_X4 U445 ( .A1(n1151), .A2(n1166), .ZN(n681) );
  XNOR2_X2 U446 ( .A(n698), .B(n546), .ZN(product[49]) );
  AOI21_X4 U458 ( .B1(n3480), .B2(n703), .A(n695), .ZN(n693) );
  NAND2_X4 U461 ( .A1(n992), .A2(n697), .ZN(n546) );
  NOR2_X4 U463 ( .A1(n1167), .A2(n1182), .ZN(n696) );
  NAND2_X4 U467 ( .A1(n993), .A2(n700), .ZN(n547) );
  NAND2_X4 U470 ( .A1(n1183), .A2(n1200), .ZN(n700) );
  XNOR2_X2 U479 ( .A(n717), .B(n549), .ZN(product[46]) );
  NAND2_X4 U481 ( .A1(n725), .A2(n709), .ZN(n707) );
  AOI21_X4 U482 ( .B1(n726), .B2(n709), .A(n710), .ZN(n708) );
  NAND2_X4 U533 ( .A1(n999), .A2(n748), .ZN(n553) );
  XOR2_X2 U537 ( .A(n756), .B(n554), .Z(product[41]) );
  NAND2_X4 U543 ( .A1(n1000), .A2(n755), .ZN(n554) );
  NAND2_X4 U551 ( .A1(n757), .A2(n760), .ZN(n555) );
  AOI21_X4 U557 ( .B1(n806), .B2(n763), .A(n764), .ZN(n531) );
  NAND2_X4 U570 ( .A1(n1003), .A2(n773), .ZN(n557) );
  XNOR2_X2 U574 ( .A(n779), .B(n558), .ZN(product[37]) );
  XOR2_X2 U582 ( .A(n782), .B(n559), .Z(product[36]) );
  XOR2_X2 U588 ( .A(n790), .B(n560), .Z(product[35]) );
  XNOR2_X2 U599 ( .A(n795), .B(n561), .ZN(product[34]) );
  AOI21_X4 U600 ( .B1(n795), .B2(n791), .A(n792), .ZN(n790) );
  XNOR2_X2 U607 ( .A(n802), .B(n562), .ZN(product[33]) );
  OAI21_X4 U608 ( .B1(n805), .B2(n796), .A(n797), .ZN(n795) );
  XOR2_X2 U617 ( .A(n805), .B(n563), .Z(product[32]) );
  XNOR2_X2 U623 ( .A(n813), .B(n564), .ZN(product[31]) );
  XOR2_X2 U634 ( .A(n816), .B(n565), .Z(product[30]) );
  XOR2_X2 U640 ( .A(n821), .B(n566), .Z(product[29]) );
  NAND2_X4 U644 ( .A1(n1012), .A2(n820), .ZN(n566) );
  XNOR2_X2 U648 ( .A(n826), .B(n567), .ZN(product[28]) );
  AOI21_X4 U649 ( .B1(n826), .B2(n822), .A(n823), .ZN(n821) );
  XOR2_X2 U656 ( .A(n836), .B(n568), .Z(product[27]) );
  NOR2_X4 U659 ( .A1(n830), .A2(n842), .ZN(n828) );
  NAND2_X4 U665 ( .A1(n3514), .A2(n835), .ZN(n568) );
  XNOR2_X2 U669 ( .A(n841), .B(n569), .ZN(product[26]) );
  XNOR2_X2 U677 ( .A(n848), .B(n570), .ZN(product[25]) );
  XOR2_X2 U687 ( .A(n855), .B(n571), .Z(product[24]) );
  XOR2_X2 U708 ( .A(n866), .B(n573), .Z(product[22]) );
  OAI21_X4 U709 ( .B1(n866), .B2(n864), .A(n865), .ZN(n863) );
  NAND2_X4 U710 ( .A1(n1019), .A2(n865), .ZN(n573) );
  XOR2_X2 U714 ( .A(n871), .B(n574), .Z(product[21]) );
  AOI21_X4 U715 ( .B1(n876), .B2(n867), .A(n868), .ZN(n866) );
  NOR2_X4 U716 ( .A1(n869), .A2(n874), .ZN(n867) );
  OAI21_X4 U717 ( .B1(n869), .B2(n875), .A(n870), .ZN(n868) );
  NAND2_X4 U718 ( .A1(n1020), .A2(n870), .ZN(n574) );
  NOR2_X4 U720 ( .A1(n1862), .A2(n1881), .ZN(n869) );
  NAND2_X4 U721 ( .A1(n1862), .A2(n1881), .ZN(n870) );
  XNOR2_X2 U722 ( .A(n876), .B(n575), .ZN(product[20]) );
  AOI21_X4 U723 ( .B1(n876), .B2(n872), .A(n873), .ZN(n871) );
  NAND2_X4 U726 ( .A1(n872), .A2(n875), .ZN(n575) );
  XNOR2_X2 U730 ( .A(n882), .B(n576), .ZN(product[19]) );
  NOR2_X4 U733 ( .A1(n883), .A2(n880), .ZN(n878) );
  NAND2_X4 U735 ( .A1(n1022), .A2(n881), .ZN(n576) );
  NOR2_X4 U737 ( .A1(n1900), .A2(n1917), .ZN(n880) );
  NAND2_X4 U738 ( .A1(n1900), .A2(n1917), .ZN(n881) );
  XNOR2_X2 U739 ( .A(n889), .B(n577), .ZN(product[18]) );
  XOR2_X2 U749 ( .A(n896), .B(n578), .Z(product[17]) );
  OAI21_X4 U750 ( .B1(n896), .B2(n890), .A(n891), .ZN(n889) );
  NAND2_X4 U755 ( .A1(n892), .A2(n891), .ZN(n578) );
  XOR2_X2 U759 ( .A(n904), .B(n579), .Z(product[16]) );
  OAI21_X4 U761 ( .B1(n898), .B2(n915), .A(n899), .ZN(n897) );
  NAND2_X4 U762 ( .A1(n905), .A2(n900), .ZN(n898) );
  AOI21_X4 U763 ( .B1(n906), .B2(n900), .A(n901), .ZN(n899) );
  NAND2_X4 U766 ( .A1(n900), .A2(n903), .ZN(n579) );
  XOR2_X2 U770 ( .A(n909), .B(n580), .Z(product[15]) );
  AOI21_X4 U771 ( .B1(n914), .B2(n905), .A(n906), .ZN(n904) );
  NOR2_X4 U772 ( .A1(n907), .A2(n912), .ZN(n905) );
  OAI21_X4 U773 ( .B1(n907), .B2(n913), .A(n908), .ZN(n906) );
  NAND2_X4 U774 ( .A1(n1026), .A2(n908), .ZN(n580) );
  NOR2_X4 U776 ( .A1(n1964), .A2(n1977), .ZN(n907) );
  NAND2_X4 U777 ( .A1(n1964), .A2(n1977), .ZN(n908) );
  XNOR2_X2 U778 ( .A(n914), .B(n581), .ZN(product[14]) );
  AOI21_X4 U779 ( .B1(n914), .B2(n910), .A(n911), .ZN(n909) );
  NAND2_X4 U782 ( .A1(n910), .A2(n913), .ZN(n581) );
  NOR2_X4 U784 ( .A1(n1978), .A2(n1989), .ZN(n912) );
  NAND2_X4 U785 ( .A1(n1978), .A2(n1989), .ZN(n913) );
  XNOR2_X2 U786 ( .A(n920), .B(n582), .ZN(product[13]) );
  AOI21_X4 U788 ( .B1(n916), .B2(n924), .A(n917), .ZN(n915) );
  NOR2_X4 U789 ( .A1(n918), .A2(n921), .ZN(n916) );
  OAI21_X4 U790 ( .B1(n918), .B2(n922), .A(n919), .ZN(n917) );
  NAND2_X4 U791 ( .A1(n1028), .A2(n919), .ZN(n582) );
  NOR2_X4 U793 ( .A1(n1990), .A2(n2001), .ZN(n918) );
  NAND2_X4 U794 ( .A1(n1990), .A2(n2001), .ZN(n919) );
  XOR2_X2 U795 ( .A(n923), .B(n583), .Z(product[12]) );
  OAI21_X4 U796 ( .B1(n923), .B2(n921), .A(n922), .ZN(n920) );
  NAND2_X4 U797 ( .A1(n1029), .A2(n922), .ZN(n583) );
  NOR2_X4 U799 ( .A1(n2002), .A2(n2011), .ZN(n921) );
  NAND2_X4 U800 ( .A1(n2002), .A2(n2011), .ZN(n922) );
  XOR2_X2 U801 ( .A(n931), .B(n584), .Z(product[11]) );
  OAI21_X4 U803 ( .B1(n925), .B2(n937), .A(n926), .ZN(n924) );
  NAND2_X4 U804 ( .A1(n932), .A2(n927), .ZN(n925) );
  AOI21_X4 U805 ( .B1(n927), .B2(n933), .A(n928), .ZN(n926) );
  NAND2_X4 U808 ( .A1(n927), .A2(n930), .ZN(n584) );
  NOR2_X4 U810 ( .A1(n2012), .A2(n2021), .ZN(n929) );
  NAND2_X4 U811 ( .A1(n2012), .A2(n2021), .ZN(n930) );
  XNOR2_X2 U812 ( .A(n585), .B(n936), .ZN(product[10]) );
  AOI21_X4 U813 ( .B1(n936), .B2(n932), .A(n933), .ZN(n931) );
  NAND2_X4 U816 ( .A1(n932), .A2(n935), .ZN(n585) );
  XNOR2_X2 U820 ( .A(n586), .B(n942), .ZN(product[9]) );
  AOI21_X4 U822 ( .B1(n942), .B2(n938), .A(n939), .ZN(n937) );
  NAND2_X4 U825 ( .A1(n938), .A2(n941), .ZN(n586) );
  NOR2_X4 U827 ( .A1(n2030), .A2(n2037), .ZN(n940) );
  NAND2_X4 U828 ( .A1(n2030), .A2(n2037), .ZN(n941) );
  XOR2_X2 U829 ( .A(n949), .B(n587), .Z(product[8]) );
  OAI21_X4 U830 ( .B1(n943), .B2(n955), .A(n944), .ZN(n942) );
  NAND2_X4 U831 ( .A1(n945), .A2(n950), .ZN(n943) );
  AOI21_X4 U832 ( .B1(n945), .B2(n951), .A(n946), .ZN(n944) );
  NAND2_X4 U835 ( .A1(n945), .A2(n948), .ZN(n587) );
  NOR2_X4 U837 ( .A1(n2038), .A2(n2043), .ZN(n947) );
  NAND2_X4 U838 ( .A1(n2038), .A2(n2043), .ZN(n948) );
  XNOR2_X2 U839 ( .A(n954), .B(n588), .ZN(product[7]) );
  AOI21_X4 U840 ( .B1(n954), .B2(n950), .A(n951), .ZN(n949) );
  NAND2_X4 U843 ( .A1(n950), .A2(n953), .ZN(n588) );
  NOR2_X4 U845 ( .A1(n2044), .A2(n2049), .ZN(n952) );
  NAND2_X4 U846 ( .A1(n2044), .A2(n2049), .ZN(n953) );
  XNOR2_X2 U847 ( .A(n589), .B(n960), .ZN(product[6]) );
  AOI21_X4 U849 ( .B1(n956), .B2(n960), .A(n957), .ZN(n955) );
  NAND2_X4 U852 ( .A1(n956), .A2(n959), .ZN(n589) );
  NOR2_X4 U854 ( .A1(n2050), .A2(n2053), .ZN(n958) );
  NAND2_X4 U855 ( .A1(n2050), .A2(n2053), .ZN(n959) );
  XOR2_X2 U856 ( .A(n590), .B(n963), .Z(product[5]) );
  OAI21_X4 U857 ( .B1(n961), .B2(n963), .A(n962), .ZN(n960) );
  NAND2_X4 U858 ( .A1(n1036), .A2(n962), .ZN(n590) );
  NOR2_X4 U860 ( .A1(n2054), .A2(n2057), .ZN(n961) );
  NAND2_X4 U861 ( .A1(n2054), .A2(n2057), .ZN(n962) );
  XNOR2_X2 U862 ( .A(n591), .B(n968), .ZN(product[4]) );
  AOI21_X4 U863 ( .B1(n964), .B2(n968), .A(n965), .ZN(n963) );
  NAND2_X4 U866 ( .A1(n964), .A2(n967), .ZN(n591) );
  NOR2_X4 U868 ( .A1(n2058), .A2(n2059), .ZN(n966) );
  NAND2_X4 U869 ( .A1(n2058), .A2(n2059), .ZN(n967) );
  XOR2_X2 U870 ( .A(n592), .B(n971), .Z(product[3]) );
  OAI21_X4 U871 ( .B1(n969), .B2(n971), .A(n970), .ZN(n968) );
  NAND2_X4 U872 ( .A1(n1038), .A2(n970), .ZN(n592) );
  NOR2_X4 U874 ( .A1(n2060), .A2(n2075), .ZN(n969) );
  NAND2_X4 U875 ( .A1(n2060), .A2(n2075), .ZN(n970) );
  XNOR2_X2 U876 ( .A(n593), .B(n976), .ZN(product[2]) );
  AOI21_X4 U877 ( .B1(n972), .B2(n976), .A(n973), .ZN(n971) );
  NAND2_X4 U880 ( .A1(n972), .A2(n975), .ZN(n593) );
  NOR2_X4 U882 ( .A1(n2603), .A2(n2635), .ZN(n974) );
  NAND2_X4 U883 ( .A1(n2603), .A2(n2635), .ZN(n975) );
  NAND2_X4 U886 ( .A1(n1040), .A2(n978), .ZN(n594) );
  NOR2_X4 U888 ( .A1(n2636), .A2(n2076), .ZN(n977) );
  NAND2_X4 U889 ( .A1(n2636), .A2(n2076), .ZN(n978) );
  FA_X1 U890 ( .A(n2095), .B(n1045), .CI(n1048), .CO(n1042), .S(n1043) );
  FA_X1 U892 ( .A(n1052), .B(n2128), .CI(n1049), .CO(n1046), .S(n1047) );
  FA_X1 U893 ( .A(n2078), .B(n1054), .CI(n2096), .CO(n1048), .S(n1049) );
  FA_X1 U894 ( .A(n1053), .B(n1060), .CI(n1058), .CO(n1050), .S(n1051) );
  FA_X1 U895 ( .A(n2129), .B(n1055), .CI(n2097), .CO(n1052), .S(n1053) );
  FA_X1 U897 ( .A(n1064), .B(n1061), .CI(n1059), .CO(n1056), .S(n1057) );
  FA_X1 U898 ( .A(n2162), .B(n2098), .CI(n1066), .CO(n1058), .S(n1059) );
  FA_X1 U899 ( .A(n2079), .B(n1068), .CI(n2130), .CO(n1060), .S(n1061) );
  FA_X1 U900 ( .A(n1072), .B(n1067), .CI(n1065), .CO(n1062), .S(n1063) );
  FA_X1 U901 ( .A(n1076), .B(n2099), .CI(n1074), .CO(n1064), .S(n1065) );
  FA_X1 U902 ( .A(n2163), .B(n1069), .CI(n2131), .CO(n1066), .S(n1067) );
  FA_X1 U904 ( .A(n1080), .B(n1082), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U905 ( .A(n1077), .B(n1084), .CI(n1075), .CO(n1072), .S(n1073) );
  FA_X1 U906 ( .A(n2132), .B(n2100), .CI(n2196), .CO(n1074), .S(n1075) );
  FA_X1 U907 ( .A(n2080), .B(n1086), .CI(n2164), .CO(n1076), .S(n1077) );
  FA_X1 U908 ( .A(n1090), .B(n1083), .CI(n1081), .CO(n1078), .S(n1079) );
  FA_X1 U909 ( .A(n1085), .B(n1094), .CI(n1092), .CO(n1080), .S(n1081) );
  FA_X1 U910 ( .A(n2101), .B(n2133), .CI(n1096), .CO(n1082), .S(n1083) );
  FA_X1 U911 ( .A(n2197), .B(n1087), .CI(n2165), .CO(n1084), .S(n1085) );
  FA_X1 U913 ( .A(n1100), .B(n1093), .CI(n1091), .CO(n1088), .S(n1089) );
  FA_X1 U914 ( .A(n1095), .B(n1097), .CI(n1102), .CO(n1090), .S(n1091) );
  FA_X1 U915 ( .A(n1106), .B(n2230), .CI(n1104), .CO(n1092), .S(n1093) );
  FA_X1 U916 ( .A(n2102), .B(n2134), .CI(n2198), .CO(n1094), .S(n1095) );
  FA_X1 U917 ( .A(n2081), .B(n1108), .CI(n2166), .CO(n1096), .S(n1097) );
  FA_X1 U918 ( .A(n1112), .B(n1103), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U919 ( .A(n1116), .B(n1105), .CI(n1114), .CO(n1100), .S(n1101) );
  FA_X1 U920 ( .A(n1118), .B(n1120), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U921 ( .A(n2135), .B(n2103), .CI(n2167), .CO(n1104), .S(n1105) );
  FA_X1 U922 ( .A(n2231), .B(n1109), .CI(n2199), .CO(n1106), .S(n1107) );
  FA_X1 U924 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U925 ( .A(n1117), .B(n1128), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U926 ( .A(n1121), .B(n1130), .CI(n1119), .CO(n1114), .S(n1115) );
  FA_X1 U927 ( .A(n2264), .B(n2136), .CI(n1132), .CO(n1116), .S(n1117) );
  FA_X1 U928 ( .A(n2104), .B(n2168), .CI(n2232), .CO(n1118), .S(n1119) );
  FA_X1 U929 ( .A(n2082), .B(n1134), .CI(n2200), .CO(n1120), .S(n1121) );
  FA_X1 U930 ( .A(n1138), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U931 ( .A(n1129), .B(n1142), .CI(n1140), .CO(n1124), .S(n1125) );
  FA_X1 U932 ( .A(n1133), .B(n1144), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U933 ( .A(n1148), .B(n2137), .CI(n1146), .CO(n1128), .S(n1129) );
  FA_X1 U934 ( .A(n2105), .B(n2201), .CI(n2169), .CO(n1130), .S(n1131) );
  FA_X1 U935 ( .A(n2265), .B(n1135), .CI(n2233), .CO(n1132), .S(n1133) );
  FA_X1 U937 ( .A(n1152), .B(n1141), .CI(n1139), .CO(n1136), .S(n1137) );
  FA_X1 U938 ( .A(n1143), .B(n1156), .CI(n1154), .CO(n1138), .S(n1139) );
  FA_X1 U939 ( .A(n1145), .B(n1147), .CI(n1158), .CO(n1140), .S(n1141) );
  FA_X1 U940 ( .A(n1160), .B(n1162), .CI(n1149), .CO(n1142), .S(n1143) );
  FA_X1 U941 ( .A(n2266), .B(n2106), .CI(n2298), .CO(n1144), .S(n1145) );
  FA_X1 U942 ( .A(n2138), .B(n2170), .CI(n2234), .CO(n1146), .S(n1147) );
  FA_X1 U943 ( .A(n2083), .B(n1164), .CI(n2202), .CO(n1148), .S(n1149) );
  FA_X1 U944 ( .A(n1168), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U945 ( .A(n1157), .B(n1172), .CI(n1170), .CO(n1152), .S(n1153) );
  FA_X1 U946 ( .A(n1174), .B(n1161), .CI(n1159), .CO(n1154), .S(n1155) );
  FA_X1 U947 ( .A(n1176), .B(n1178), .CI(n1163), .CO(n1156), .S(n1157) );
  FA_X1 U948 ( .A(n2171), .B(n2203), .CI(n1180), .CO(n1158), .S(n1159) );
  FA_X1 U949 ( .A(n2107), .B(n2235), .CI(n2139), .CO(n1160), .S(n1161) );
  FA_X1 U950 ( .A(n2299), .B(n1165), .CI(n2267), .CO(n1162), .S(n1163) );
  FA_X1 U952 ( .A(n1184), .B(n1171), .CI(n1169), .CO(n1166), .S(n1167) );
  FA_X1 U953 ( .A(n1173), .B(n1188), .CI(n1186), .CO(n1168), .S(n1169) );
  FA_X1 U954 ( .A(n1190), .B(n1179), .CI(n1175), .CO(n1170), .S(n1171) );
  FA_X1 U955 ( .A(n1181), .B(n1192), .CI(n1177), .CO(n1172), .S(n1173) );
  FA_X1 U956 ( .A(n1196), .B(n2332), .CI(n1194), .CO(n1174), .S(n1175) );
  FA_X1 U957 ( .A(n2268), .B(n2140), .CI(n2300), .CO(n1176), .S(n1177) );
  FA_X1 U958 ( .A(n2108), .B(n2204), .CI(n2172), .CO(n1178), .S(n1179) );
  FA_X1 U959 ( .A(n2084), .B(n1198), .CI(n2236), .CO(n1180), .S(n1181) );
  FA_X1 U960 ( .A(n1202), .B(n1187), .CI(n1185), .CO(n1182), .S(n1183) );
  FA_X1 U961 ( .A(n1189), .B(n1206), .CI(n1204), .CO(n1184), .S(n1185) );
  FA_X1 U962 ( .A(n1208), .B(n1210), .CI(n1191), .CO(n1186), .S(n1187) );
  FA_X1 U963 ( .A(n1193), .B(n1197), .CI(n1195), .CO(n1188), .S(n1189) );
  FA_X1 U964 ( .A(n1214), .B(n1216), .CI(n1212), .CO(n1190), .S(n1191) );
  FA_X1 U965 ( .A(n2141), .B(n2205), .CI(n2173), .CO(n1192), .S(n1193) );
  FA_X1 U966 ( .A(n2109), .B(n2269), .CI(n2237), .CO(n1194), .S(n1195) );
  FA_X1 U967 ( .A(n2333), .B(n1199), .CI(n2301), .CO(n1196), .S(n1197) );
  FA_X1 U969 ( .A(n1220), .B(n1205), .CI(n1203), .CO(n1200), .S(n1201) );
  FA_X1 U970 ( .A(n1207), .B(n1224), .CI(n1222), .CO(n1202), .S(n1203) );
  FA_X1 U971 ( .A(n1211), .B(n1226), .CI(n1209), .CO(n1204), .S(n1205) );
  FA_X1 U972 ( .A(n1215), .B(n1213), .CI(n1228), .CO(n1206), .S(n1207) );
  FA_X1 U973 ( .A(n1230), .B(n1232), .CI(n1217), .CO(n1208), .S(n1209) );
  FA_X1 U974 ( .A(n2366), .B(n2334), .CI(n1234), .CO(n1210), .S(n1211) );
  FA_X1 U975 ( .A(n2302), .B(n2174), .CI(n2270), .CO(n1212), .S(n1213) );
  FA_X1 U976 ( .A(n2142), .B(n2206), .CI(n2110), .CO(n1214), .S(n1215) );
  FA_X1 U977 ( .A(n2085), .B(n1236), .CI(n2238), .CO(n1216), .S(n1217) );
  FA_X1 U978 ( .A(n1240), .B(n1223), .CI(n1221), .CO(n1218), .S(n1219) );
  FA_X1 U979 ( .A(n1225), .B(n1244), .CI(n1242), .CO(n1220), .S(n1221) );
  FA_X1 U980 ( .A(n1246), .B(n1229), .CI(n1227), .CO(n1222), .S(n1223) );
  FA_X1 U981 ( .A(n1233), .B(n1231), .CI(n1248), .CO(n1224), .S(n1225) );
  FA_X1 U982 ( .A(n1250), .B(n1252), .CI(n1235), .CO(n1226), .S(n1227) );
  FA_X1 U983 ( .A(n1256), .B(n2239), .CI(n1254), .CO(n1228), .S(n1229) );
  FA_X1 U984 ( .A(n2175), .B(n2271), .CI(n2207), .CO(n1230), .S(n1231) );
  FA_X1 U985 ( .A(n2111), .B(n2303), .CI(n2143), .CO(n1232), .S(n1233) );
  FA_X1 U986 ( .A(n2367), .B(n1237), .CI(n2335), .CO(n1234), .S(n1235) );
  FA_X1 U988 ( .A(n1260), .B(n1243), .CI(n1241), .CO(n1238), .S(n1239) );
  FA_X1 U989 ( .A(n1245), .B(n1264), .CI(n1262), .CO(n1240), .S(n1241) );
  FA_X1 U990 ( .A(n1249), .B(n1266), .CI(n1247), .CO(n1242), .S(n1243) );
  FA_X1 U991 ( .A(n1270), .B(n1251), .CI(n1268), .CO(n1244), .S(n1245) );
  FA_X1 U992 ( .A(n1253), .B(n1257), .CI(n1255), .CO(n1246), .S(n1247) );
  FA_X1 U993 ( .A(n1272), .B(n1276), .CI(n1274), .CO(n1248), .S(n1249) );
  FA_X1 U994 ( .A(n2336), .B(n2368), .CI(n2400), .CO(n1250), .S(n1251) );
  FA_X1 U995 ( .A(n2304), .B(n2144), .CI(n2208), .CO(n1252), .S(n1253) );
  FA_X1 U996 ( .A(n2112), .B(n2240), .CI(n2176), .CO(n1254), .S(n1255) );
  FA_X1 U997 ( .A(n2086), .B(n1278), .CI(n2272), .CO(n1256), .S(n1257) );
  FA_X1 U998 ( .A(n1282), .B(n1263), .CI(n1261), .CO(n1258), .S(n1259) );
  FA_X1 U999 ( .A(n1265), .B(n1286), .CI(n1284), .CO(n1260), .S(n1261) );
  FA_X1 U1000 ( .A(n1269), .B(n1288), .CI(n1267), .CO(n1262), .S(n1263) );
  FA_X1 U1001 ( .A(n1271), .B(n1292), .CI(n1290), .CO(n1264), .S(n1265) );
  FA_X1 U1002 ( .A(n1273), .B(n1277), .CI(n1275), .CO(n1266), .S(n1267) );
  FA_X1 U1003 ( .A(n1294), .B(n1298), .CI(n1296), .CO(n1268), .S(n1269) );
  FA_X1 U1004 ( .A(n2273), .B(n2305), .CI(n1300), .CO(n1270), .S(n1271) );
  FA_X1 U1005 ( .A(n2177), .B(n2241), .CI(n2209), .CO(n1272), .S(n1273) );
  FA_X1 U1006 ( .A(n2113), .B(n2337), .CI(n2145), .CO(n1274), .S(n1275) );
  FA_X1 U1007 ( .A(n2401), .B(n1279), .CI(n2369), .CO(n1276), .S(n1277) );
  FA_X1 U1009 ( .A(n1285), .B(n1304), .CI(n1283), .CO(n1280), .S(n1281) );
  FA_X1 U1010 ( .A(n1287), .B(n1308), .CI(n1306), .CO(n1282), .S(n1283) );
  FA_X1 U1011 ( .A(n1310), .B(n1291), .CI(n1289), .CO(n1284), .S(n1285) );
  FA_X1 U1012 ( .A(n1293), .B(n1314), .CI(n1312), .CO(n1286), .S(n1287) );
  FA_X1 U1013 ( .A(n1295), .B(n1297), .CI(n1299), .CO(n1288), .S(n1289) );
  FA_X1 U1014 ( .A(n1316), .B(n1318), .CI(n1301), .CO(n1290), .S(n1291) );
  FA_X1 U1015 ( .A(n1322), .B(n2434), .CI(n1320), .CO(n1292), .S(n1293) );
  FA_X1 U1016 ( .A(n2210), .B(n2402), .CI(n2370), .CO(n1294), .S(n1295) );
  FA_X1 U1017 ( .A(n2178), .B(n2306), .CI(n2338), .CO(n1296), .S(n1297) );
  FA_X1 U1018 ( .A(n2114), .B(n2146), .CI(n2242), .CO(n1298), .S(n1299) );
  FA_X1 U1019 ( .A(n2087), .B(n1324), .CI(n2274), .CO(n1300), .S(n1301) );
  FA_X1 U1020 ( .A(n1328), .B(n1307), .CI(n1305), .CO(n1302), .S(n1303) );
  FA_X1 U1021 ( .A(n1309), .B(n1332), .CI(n1330), .CO(n1304), .S(n1305) );
  FA_X1 U1022 ( .A(n1334), .B(n1313), .CI(n1311), .CO(n1306), .S(n1307) );
  FA_X1 U1023 ( .A(n1315), .B(n1338), .CI(n1336), .CO(n1308), .S(n1309) );
  FA_X1 U1024 ( .A(n1321), .B(n1319), .CI(n1340), .CO(n1310), .S(n1311) );
  FA_X1 U1025 ( .A(n1323), .B(n1342), .CI(n1317), .CO(n1312), .S(n1313) );
  FA_X1 U1026 ( .A(n1346), .B(n1348), .CI(n1344), .CO(n1314), .S(n1315) );
  FA_X1 U1027 ( .A(n2275), .B(n2307), .CI(n2243), .CO(n1316), .S(n1317) );
  FA_X1 U1028 ( .A(n2339), .B(n2179), .CI(n2211), .CO(n1318), .S(n1319) );
  FA_X1 U1029 ( .A(n2115), .B(n2371), .CI(n2147), .CO(n1320), .S(n1321) );
  FA_X1 U1030 ( .A(n2435), .B(n1325), .CI(n2403), .CO(n1322), .S(n1323) );
  FA_X1 U1032 ( .A(n1352), .B(n1331), .CI(n1329), .CO(n1326), .S(n1327) );
  FA_X1 U1033 ( .A(n1333), .B(n1356), .CI(n1354), .CO(n1328), .S(n1329) );
  FA_X1 U1034 ( .A(n1358), .B(n1337), .CI(n1335), .CO(n1330), .S(n1331) );
  FA_X1 U1035 ( .A(n1360), .B(n1341), .CI(n1339), .CO(n1332), .S(n1333) );
  FA_X1 U1036 ( .A(n1364), .B(n1347), .CI(n1362), .CO(n1334), .S(n1335) );
  FA_X1 U1037 ( .A(n1343), .B(n1349), .CI(n1345), .CO(n1336), .S(n1337) );
  FA_X1 U1038 ( .A(n1366), .B(n1370), .CI(n1368), .CO(n1338), .S(n1339) );
  FA_X1 U1039 ( .A(n2468), .B(n2436), .CI(n1372), .CO(n1340), .S(n1341) );
  FA_X1 U1040 ( .A(n2212), .B(n2404), .CI(n2372), .CO(n1342), .S(n1343) );
  FA_X1 U1041 ( .A(n2116), .B(n2340), .CI(n2244), .CO(n1344), .S(n1345) );
  FA_X1 U1042 ( .A(n2148), .B(n2276), .CI(n2180), .CO(n1346), .S(n1347) );
  FA_X1 U1043 ( .A(n2088), .B(n1374), .CI(n2308), .CO(n1348), .S(n1349) );
  FA_X1 U1045 ( .A(n1357), .B(n1382), .CI(n1380), .CO(n1352), .S(n1353) );
  FA_X1 U1047 ( .A(n1386), .B(n1365), .CI(n1363), .CO(n1356), .S(n1357) );
  FA_X1 U1048 ( .A(n1390), .B(n1369), .CI(n1388), .CO(n1358), .S(n1359) );
  FA_X1 U1049 ( .A(n1367), .B(n1373), .CI(n1371), .CO(n1360), .S(n1361) );
  FA_X1 U1050 ( .A(n1394), .B(n1396), .CI(n1392), .CO(n1362), .S(n1363) );
  FA_X1 U1051 ( .A(n1400), .B(n2341), .CI(n1398), .CO(n1364), .S(n1365) );
  FA_X1 U1052 ( .A(n2309), .B(n2373), .CI(n2245), .CO(n1366), .S(n1367) );
  FA_X1 U1053 ( .A(n2181), .B(n2405), .CI(n2213), .CO(n1368), .S(n1369) );
  FA_X1 U1054 ( .A(n2117), .B(n2437), .CI(n2149), .CO(n1370), .S(n1371) );
  FA_X1 U1055 ( .A(n2469), .B(n1375), .CI(n2277), .CO(n1372), .S(n1373) );
  FA_X1 U1059 ( .A(n1410), .B(n1387), .CI(n1385), .CO(n1380), .S(n1381) );
  FA_X1 U1060 ( .A(n1389), .B(n1391), .CI(n1412), .CO(n1382), .S(n1383) );
  FA_X1 U1061 ( .A(n1416), .B(n1418), .CI(n1414), .CO(n1384), .S(n1385) );
  FA_X1 U1062 ( .A(n1399), .B(n1397), .CI(n1393), .CO(n1386), .S(n1387) );
  FA_X1 U1063 ( .A(n1401), .B(n1422), .CI(n1395), .CO(n1388), .S(n1389) );
  FA_X1 U1064 ( .A(n1420), .B(n1426), .CI(n1424), .CO(n1390), .S(n1391) );
  FA_X1 U1065 ( .A(n2438), .B(n2470), .CI(n2502), .CO(n1392), .S(n1393) );
  FA_X1 U1066 ( .A(n2406), .B(n2374), .CI(n2246), .CO(n1394), .S(n1395) );
  FA_X1 U1067 ( .A(n2214), .B(n2310), .CI(n2118), .CO(n1396), .S(n1397) );
  FA_X1 U1068 ( .A(n2150), .B(n2182), .CI(n2278), .CO(n1398), .S(n1399) );
  FA_X1 U1069 ( .A(n2089), .B(n1428), .CI(n2342), .CO(n1400), .S(n1401) );
  FA_X1 U1071 ( .A(n1409), .B(n1436), .CI(n1434), .CO(n1404), .S(n1405) );
  FA_X1 U1072 ( .A(n1438), .B(n1413), .CI(n1411), .CO(n1406), .S(n1407) );
  FA_X1 U1073 ( .A(n1415), .B(n1417), .CI(n1440), .CO(n1408), .S(n1409) );
  FA_X1 U1074 ( .A(n1419), .B(n1444), .CI(n1442), .CO(n1410), .S(n1411) );
  FA_X1 U1075 ( .A(n1425), .B(n1423), .CI(n1446), .CO(n1412), .S(n1413) );
  FA_X1 U1076 ( .A(n1427), .B(n1452), .CI(n1421), .CO(n1414), .S(n1415) );
  FA_X1 U1077 ( .A(n1448), .B(n1454), .CI(n1450), .CO(n1416), .S(n1417) );
  FA_X1 U1078 ( .A(n2247), .B(n2311), .CI(n1456), .CO(n1418), .S(n1419) );
  FA_X1 U1079 ( .A(n2183), .B(n2343), .CI(n2215), .CO(n1420), .S(n1421) );
  FA_X1 U1080 ( .A(n2151), .B(n2375), .CI(n2407), .CO(n1422), .S(n1423) );
  FA_X1 U1081 ( .A(n2439), .B(n2279), .CI(n2119), .CO(n1424), .S(n1425) );
  FA_X1 U1082 ( .A(n2471), .B(n1429), .CI(n2503), .CO(n1426), .S(n1427) );
  FA_X1 U1084 ( .A(n1435), .B(n1460), .CI(n1433), .CO(n1430), .S(n1431) );
  FA_X1 U1085 ( .A(n1437), .B(n1464), .CI(n1462), .CO(n1432), .S(n1433) );
  FA_X1 U1087 ( .A(n1443), .B(n1445), .CI(n1468), .CO(n1436), .S(n1437) );
  FA_X1 U1089 ( .A(n1453), .B(n1455), .CI(n1474), .CO(n1440), .S(n1441) );
  FA_X1 U1091 ( .A(n1480), .B(n1478), .CI(n1482), .CO(n1444), .S(n1445) );
  FA_X1 U1092 ( .A(n1484), .B(n2536), .CI(n1476), .CO(n1446), .S(n1447) );
  FA_X1 U1093 ( .A(n2504), .B(n2472), .CI(n2280), .CO(n1448), .S(n1449) );
  FA_X1 U1095 ( .A(n2152), .B(n2376), .CI(n2216), .CO(n1452), .S(n1453) );
  FA_X1 U1096 ( .A(n2184), .B(n2312), .CI(n2120), .CO(n1454), .S(n1455) );
  FA_X1 U1097 ( .A(n2090), .B(n1486), .CI(n2344), .CO(n1456), .S(n1457) );
  FA_X1 U1098 ( .A(n1463), .B(n1490), .CI(n1461), .CO(n1458), .S(n1459) );
  FA_X1 U1099 ( .A(n1465), .B(n1494), .CI(n1492), .CO(n1460), .S(n1461) );
  FA_X1 U1100 ( .A(n1496), .B(n1469), .CI(n1467), .CO(n1462), .S(n1463) );
  FA_X1 U1101 ( .A(n1471), .B(n1473), .CI(n1498), .CO(n1464), .S(n1465) );
  FA_X1 U1102 ( .A(n1502), .B(n1500), .CI(n1475), .CO(n1466), .S(n1467) );
  FA_X1 U1103 ( .A(n1506), .B(n1481), .CI(n1504), .CO(n1468), .S(n1469) );
  FA_X1 U1104 ( .A(n1483), .B(n1477), .CI(n1479), .CO(n1470), .S(n1471) );
  FA_X1 U1105 ( .A(n1514), .B(n1512), .CI(n1485), .CO(n1472), .S(n1473) );
  FA_X1 U1106 ( .A(n1508), .B(n1516), .CI(n1510), .CO(n1474), .S(n1475) );
  FA_X1 U1108 ( .A(n2185), .B(n2377), .CI(n2217), .CO(n1478), .S(n1479) );
  FA_X1 U1109 ( .A(n2153), .B(n2441), .CI(n2409), .CO(n1480), .S(n1481) );
  FA_X1 U1110 ( .A(n2473), .B(n2281), .CI(n2121), .CO(n1482), .S(n1483) );
  FA_X1 U1111 ( .A(n2537), .B(n1487), .CI(n2505), .CO(n1484), .S(n1485) );
  FA_X1 U1114 ( .A(n1495), .B(n1524), .CI(n1522), .CO(n1490), .S(n1491) );
  FA_X1 U1115 ( .A(n1499), .B(n1526), .CI(n1497), .CO(n1492), .S(n1493) );
  FA_X1 U1117 ( .A(n1532), .B(n1530), .CI(n1505), .CO(n1496), .S(n1497) );
  FA_X1 U1118 ( .A(n1534), .B(n1536), .CI(n1507), .CO(n1498), .S(n1499) );
  FA_X1 U1121 ( .A(n1542), .B(n1538), .CI(n1544), .CO(n1504), .S(n1505) );
  FA_X1 U1122 ( .A(n2570), .B(n2474), .CI(n1546), .CO(n1506), .S(n1507) );
  FA_X1 U1123 ( .A(n2538), .B(n2506), .CI(n2442), .CO(n1508), .S(n1509) );
  FA_X1 U1124 ( .A(n2346), .B(n2282), .CI(n2250), .CO(n1510), .S(n1511) );
  FA_X1 U1126 ( .A(n2122), .B(n2314), .CI(n2154), .CO(n1514), .S(n1515) );
  FA_X1 U1127 ( .A(n2091), .B(n1548), .CI(n2378), .CO(n1516), .S(n1517) );
  FA_X1 U1129 ( .A(n1525), .B(n1556), .CI(n1554), .CO(n1520), .S(n1521) );
  FA_X1 U1131 ( .A(n1531), .B(n1533), .CI(n1560), .CO(n1524), .S(n1525) );
  FA_X1 U1132 ( .A(n1562), .B(n1537), .CI(n1535), .CO(n1526), .S(n1527) );
  FA_X1 U1135 ( .A(n1547), .B(n1572), .CI(n1539), .CO(n1532), .S(n1533) );
  FA_X1 U1136 ( .A(n1574), .B(n1570), .CI(n1576), .CO(n1534), .S(n1535) );
  FA_X1 U1137 ( .A(n2411), .B(n2379), .CI(n1578), .CO(n1536), .S(n1537) );
  FA_X1 U1138 ( .A(n2443), .B(n2347), .CI(n2315), .CO(n1538), .S(n1539) );
  FA_X1 U1139 ( .A(n2475), .B(n2283), .CI(n2251), .CO(n1540), .S(n1541) );
  FA_X1 U1141 ( .A(n2539), .B(n2155), .CI(n2123), .CO(n1544), .S(n1545) );
  FA_X1 U1142 ( .A(n1580), .B(n2092), .CI(n2571), .CO(n1546), .S(n1547) );
  FA_X1 U1146 ( .A(n1561), .B(n1589), .CI(n1587), .CO(n1554), .S(n1555) );
  FA_X1 U1147 ( .A(n1591), .B(n1565), .CI(n1563), .CO(n1556), .S(n1557) );
  FA_X1 U1148 ( .A(n1593), .B(n1569), .CI(n1567), .CO(n1558), .S(n1559) );
  FA_X1 U1149 ( .A(n1597), .B(n1575), .CI(n1595), .CO(n1560), .S(n1561) );
  FA_X1 U1150 ( .A(n1573), .B(n1571), .CI(n1577), .CO(n1562), .S(n1563) );
  FA_X1 U1151 ( .A(n1579), .B(n1605), .CI(n1599), .CO(n1564), .S(n1565) );
  FA_X1 U1152 ( .A(n1607), .B(n1601), .CI(n1603), .CO(n1566), .S(n1567) );
  FA_X1 U1153 ( .A(n2604), .B(n2508), .CI(n1609), .CO(n1568), .S(n1569) );
  FA_X1 U1154 ( .A(n2476), .B(n2540), .CI(n2572), .CO(n1570), .S(n1571) );
  FA_X1 U1155 ( .A(n2284), .B(n2380), .CI(n2316), .CO(n1572), .S(n1573) );
  FA_X1 U1157 ( .A(n2188), .B(n2348), .CI(n2124), .CO(n1576), .S(n1577) );
  FA_X1 U1162 ( .A(n1619), .B(n1592), .CI(n1617), .CO(n1585), .S(n1586) );
  FA_X1 U1163 ( .A(n1621), .B(n1596), .CI(n1594), .CO(n1587), .S(n1588) );
  FA_X1 U1164 ( .A(n1623), .B(n1625), .CI(n1598), .CO(n1589), .S(n1590) );
  FA_X1 U1165 ( .A(n1600), .B(n1606), .CI(n1627), .CO(n1591), .S(n1592) );
  FA_X1 U1166 ( .A(n1608), .B(n1602), .CI(n1604), .CO(n1593), .S(n1594) );
  FA_X1 U1167 ( .A(n1633), .B(n1629), .CI(n1610), .CO(n1595), .S(n1596) );
  FA_X1 U1168 ( .A(n1637), .B(n1631), .CI(n1635), .CO(n1597), .S(n1598) );
  FA_X1 U1169 ( .A(n2445), .B(n2413), .CI(n1639), .CO(n1599), .S(n1600) );
  FA_X1 U1170 ( .A(n2317), .B(n2477), .CI(n2349), .CO(n1601), .S(n1602) );
  FA_X1 U1172 ( .A(n2541), .B(n2381), .CI(n2221), .CO(n1605), .S(n1606) );
  FA_X1 U1173 ( .A(n2189), .B(n2573), .CI(n2125), .CO(n1607), .S(n1608) );
  FA_X1 U1174 ( .A(n2605), .B(n2093), .CI(n2157), .CO(n1609), .S(n1610) );
  FA_X1 U1176 ( .A(n1618), .B(n1620), .CI(n1645), .CO(n1613), .S(n1614) );
  FA_X1 U1177 ( .A(n1649), .B(n1622), .CI(n1647), .CO(n1615), .S(n1616) );
  FA_X1 U1178 ( .A(n1651), .B(n1626), .CI(n1624), .CO(n1617), .S(n1618) );
  FA_X1 U1179 ( .A(n1628), .B(n1655), .CI(n1653), .CO(n1619), .S(n1620) );
  FA_X1 U1180 ( .A(n1632), .B(n1657), .CI(n1634), .CO(n1621), .S(n1622) );
  FA_X1 U1181 ( .A(n1638), .B(n1630), .CI(n1636), .CO(n1623), .S(n1624) );
  FA_X1 U1182 ( .A(n1663), .B(n1659), .CI(n1661), .CO(n1625), .S(n1626) );
  FA_X1 U1183 ( .A(n1665), .B(n1667), .CI(n1640), .CO(n1627), .S(n1628) );
  FA_X1 U1184 ( .A(n2350), .B(n2286), .CI(n2414), .CO(n1629), .S(n1630) );
  FA_X1 U1185 ( .A(n2190), .B(n2446), .CI(n2222), .CO(n1631), .S(n1632) );
  FA_X1 U1186 ( .A(n2158), .B(n2254), .CI(n2478), .CO(n1633), .S(n1634) );
  FA_X1 U1187 ( .A(n2542), .B(n2318), .CI(n2510), .CO(n1635), .S(n1636) );
  FA_X1 U1188 ( .A(n2606), .B(n2382), .CI(n2574), .CO(n1637), .S(n1638) );
  HA_X1 U1189 ( .A(n2126), .B(n2061), .CO(n1639), .S(n1640) );
  FA_X1 U1191 ( .A(n1648), .B(n1650), .CI(n1673), .CO(n1643), .S(n1644) );
  FA_X1 U1192 ( .A(n1677), .B(n1652), .CI(n1675), .CO(n1645), .S(n1646) );
  FA_X1 U1193 ( .A(n1656), .B(n1679), .CI(n1654), .CO(n1647), .S(n1648) );
  FA_X1 U1194 ( .A(n1681), .B(n1683), .CI(n1658), .CO(n1649), .S(n1650) );
  FA_X1 U1195 ( .A(n1685), .B(n1662), .CI(n1664), .CO(n1651), .S(n1652) );
  FA_X1 U1196 ( .A(n1668), .B(n1660), .CI(n1666), .CO(n1653), .S(n1654) );
  FA_X1 U1197 ( .A(n1691), .B(n1687), .CI(n1689), .CO(n1655), .S(n1656) );
  FA_X1 U1198 ( .A(n1695), .B(n2447), .CI(n1693), .CO(n1657), .S(n1658) );
  FA_X1 U1199 ( .A(n2383), .B(n2479), .CI(n2415), .CO(n1659), .S(n1660) );
  FA_X1 U1200 ( .A(n2319), .B(n2287), .CI(n2351), .CO(n1661), .S(n1662) );
  FA_X1 U1201 ( .A(n2223), .B(n2511), .CI(n2255), .CO(n1663), .S(n1664) );
  FA_X1 U1202 ( .A(n2543), .B(n2575), .CI(n2191), .CO(n1665), .S(n1666) );
  FA_X1 U1204 ( .A(n1699), .B(n1674), .CI(n1672), .CO(n1669), .S(n1670) );
  FA_X1 U1205 ( .A(n1676), .B(n1678), .CI(n1701), .CO(n1671), .S(n1672) );
  FA_X1 U1206 ( .A(n1705), .B(n1680), .CI(n1703), .CO(n1673), .S(n1674) );
  FA_X1 U1207 ( .A(n1684), .B(n1707), .CI(n1682), .CO(n1675), .S(n1676) );
  FA_X1 U1208 ( .A(n1686), .B(n1711), .CI(n1709), .CO(n1677), .S(n1678) );
  FA_X1 U1210 ( .A(n1713), .B(n1717), .CI(n1688), .CO(n1681), .S(n1682) );
  FA_X1 U1211 ( .A(n1721), .B(n1715), .CI(n1719), .CO(n1683), .S(n1684) );
  FA_X1 U1212 ( .A(n2480), .B(n2448), .CI(n1696), .CO(n1685), .S(n1686) );
  FA_X1 U1213 ( .A(n2288), .B(n2512), .CI(n2320), .CO(n1687), .S(n1688) );
  FA_X1 U1215 ( .A(n2576), .B(n2352), .CI(n2224), .CO(n1691), .S(n1692) );
  FA_X1 U1216 ( .A(n2192), .B(n2608), .CI(n2384), .CO(n1693), .S(n1694) );
  HA_X1 U1217 ( .A(n2160), .B(n2062), .CO(n1695), .S(n1696) );
  FA_X1 U1218 ( .A(n1725), .B(n1702), .CI(n1700), .CO(n1697), .S(n1698) );
  FA_X1 U1219 ( .A(n1704), .B(n1729), .CI(n1727), .CO(n1699), .S(n1700) );
  FA_X1 U1220 ( .A(n1731), .B(n1708), .CI(n1706), .CO(n1701), .S(n1702) );
  FA_X1 U1221 ( .A(n1733), .B(n1712), .CI(n1710), .CO(n1703), .S(n1704) );
  FA_X1 U1222 ( .A(n1737), .B(n1718), .CI(n1735), .CO(n1705), .S(n1706) );
  FA_X1 U1223 ( .A(n1722), .B(n1716), .CI(n1720), .CO(n1707), .S(n1708) );
  FA_X1 U1225 ( .A(n1745), .B(n1747), .CI(n1743), .CO(n1711), .S(n1712) );
  FA_X1 U1227 ( .A(n2353), .B(n2481), .CI(n2321), .CO(n1715), .S(n1716) );
  FA_X1 U1228 ( .A(n2257), .B(n2513), .CI(n2289), .CO(n1717), .S(n1718) );
  FA_X1 U1229 ( .A(n2225), .B(n2577), .CI(n2545), .CO(n1719), .S(n1720) );
  FA_X1 U1230 ( .A(n2193), .B(n2609), .CI(n2161), .CO(n1721), .S(n1722) );
  FA_X1 U1232 ( .A(n1732), .B(n1730), .CI(n1753), .CO(n1725), .S(n1726) );
  FA_X1 U1233 ( .A(n1734), .B(n1757), .CI(n1755), .CO(n1727), .S(n1728) );
  FA_X1 U1234 ( .A(n1759), .B(n1738), .CI(n1736), .CO(n1729), .S(n1730) );
  FA_X1 U1235 ( .A(n1744), .B(n1746), .CI(n1761), .CO(n1731), .S(n1732) );
  FA_X1 U1236 ( .A(n1740), .B(n1763), .CI(n1742), .CO(n1733), .S(n1734) );
  FA_X1 U1237 ( .A(n1767), .B(n1765), .CI(n1769), .CO(n1735), .S(n1736) );
  FA_X1 U1238 ( .A(n1748), .B(n2514), .CI(n1771), .CO(n1737), .S(n1738) );
  FA_X1 U1239 ( .A(n2450), .B(n2546), .CI(n2482), .CO(n1739), .S(n1740) );
  FA_X1 U1240 ( .A(n2578), .B(n2354), .CI(n2322), .CO(n1741), .S(n1742) );
  FA_X1 U1241 ( .A(n2290), .B(n2386), .CI(n2258), .CO(n1743), .S(n1744) );
  FA_X1 U1242 ( .A(n2226), .B(n2610), .CI(n2418), .CO(n1745), .S(n1746) );
  HA_X1 U1243 ( .A(n2194), .B(n2063), .CO(n1747), .S(n1748) );
  FA_X1 U1244 ( .A(n1775), .B(n1754), .CI(n1752), .CO(n1749), .S(n1750) );
  FA_X1 U1245 ( .A(n1777), .B(n1779), .CI(n1756), .CO(n1751), .S(n1752) );
  FA_X1 U1246 ( .A(n1760), .B(n1762), .CI(n1758), .CO(n1753), .S(n1754) );
  FA_X1 U1247 ( .A(n1783), .B(n1785), .CI(n1781), .CO(n1755), .S(n1756) );
  FA_X1 U1248 ( .A(n1772), .B(n1770), .CI(n1764), .CO(n1757), .S(n1758) );
  FA_X1 U1250 ( .A(n1787), .B(n1789), .CI(n1791), .CO(n1761), .S(n1762) );
  FA_X1 U1251 ( .A(n2451), .B(n2483), .CI(n1795), .CO(n1763), .S(n1764) );
  FA_X1 U1253 ( .A(n2355), .B(n2547), .CI(n2323), .CO(n1767), .S(n1768) );
  FA_X1 U1254 ( .A(n2291), .B(n2579), .CI(n2259), .CO(n1769), .S(n1770) );
  FA_X1 U1255 ( .A(n2227), .B(n2611), .CI(n2195), .CO(n1771), .S(n1772) );
  FA_X1 U1256 ( .A(n1799), .B(n1778), .CI(n1776), .CO(n1773), .S(n1774) );
  FA_X1 U1257 ( .A(n1803), .B(n1780), .CI(n1801), .CO(n1775), .S(n1776) );
  FA_X1 U1258 ( .A(n1784), .B(n1805), .CI(n1782), .CO(n1777), .S(n1778) );
  FA_X1 U1259 ( .A(n1807), .B(n1809), .CI(n1786), .CO(n1779), .S(n1780) );
  FA_X1 U1261 ( .A(n1811), .B(n1813), .CI(n1788), .CO(n1783), .S(n1784) );
  FA_X1 U1262 ( .A(n1815), .B(n1796), .CI(n1817), .CO(n1785), .S(n1786) );
  FA_X1 U1263 ( .A(n2356), .B(n2484), .CI(n2452), .CO(n1787), .S(n1788) );
  FA_X1 U1264 ( .A(n2292), .B(n2516), .CI(n2324), .CO(n1789), .S(n1790) );
  FA_X1 U1265 ( .A(n2580), .B(n2388), .CI(n2548), .CO(n1791), .S(n1792) );
  HA_X1 U1267 ( .A(n2228), .B(n2064), .CO(n1795), .S(n1796) );
  FA_X1 U1268 ( .A(n1821), .B(n1802), .CI(n1800), .CO(n1797), .S(n1798) );
  FA_X1 U1269 ( .A(n1804), .B(n1825), .CI(n1823), .CO(n1799), .S(n1800) );
  FA_X1 U1270 ( .A(n1808), .B(n1827), .CI(n1806), .CO(n1801), .S(n1802) );
  FA_X1 U1271 ( .A(n1829), .B(n1831), .CI(n1810), .CO(n1803), .S(n1804) );
  FA_X1 U1272 ( .A(n1818), .B(n1814), .CI(n1816), .CO(n1805), .S(n1806) );
  FA_X1 U1273 ( .A(n1833), .B(n1835), .CI(n1812), .CO(n1807), .S(n1808) );
  FA_X1 U1274 ( .A(n1839), .B(n2453), .CI(n1837), .CO(n1809), .S(n1810) );
  FA_X1 U1275 ( .A(n2389), .B(n2485), .CI(n2421), .CO(n1811), .S(n1812) );
  FA_X1 U1276 ( .A(n2357), .B(n2549), .CI(n2517), .CO(n1813), .S(n1814) );
  FA_X1 U1277 ( .A(n2325), .B(n2581), .CI(n2293), .CO(n1815), .S(n1816) );
  FA_X1 U1278 ( .A(n2229), .B(n2613), .CI(n2261), .CO(n1817), .S(n1818) );
  FA_X1 U1279 ( .A(n1843), .B(n1824), .CI(n1822), .CO(n1819), .S(n1820) );
  FA_X1 U1280 ( .A(n1845), .B(n1828), .CI(n1826), .CO(n1821), .S(n1822) );
  FA_X1 U1281 ( .A(n1830), .B(n1849), .CI(n1847), .CO(n1823), .S(n1824) );
  FA_X1 U1282 ( .A(n1851), .B(n1838), .CI(n1832), .CO(n1825), .S(n1826) );
  FA_X1 U1283 ( .A(n1834), .B(n1857), .CI(n1836), .CO(n1827), .S(n1828) );
  FA_X1 U1284 ( .A(n1853), .B(n1859), .CI(n1855), .CO(n1829), .S(n1830) );
  FA_X1 U1285 ( .A(n2486), .B(n2518), .CI(n1840), .CO(n1831), .S(n1832) );
  FA_X1 U1286 ( .A(n2358), .B(n2550), .CI(n2390), .CO(n1833), .S(n1834) );
  FA_X1 U1287 ( .A(n2582), .B(n2422), .CI(n2326), .CO(n1835), .S(n1836) );
  FA_X1 U1288 ( .A(n2614), .B(n2454), .CI(n2294), .CO(n1837), .S(n1838) );
  HA_X1 U1289 ( .A(n2262), .B(n2065), .CO(n1839), .S(n1840) );
  FA_X1 U1290 ( .A(n1863), .B(n1846), .CI(n1844), .CO(n1841), .S(n1842) );
  FA_X1 U1291 ( .A(n1848), .B(n1850), .CI(n1865), .CO(n1843), .S(n1844) );
  FA_X1 U1292 ( .A(n1852), .B(n1869), .CI(n1867), .CO(n1845), .S(n1846) );
  FA_X1 U1293 ( .A(n1860), .B(n1858), .CI(n1871), .CO(n1847), .S(n1848) );
  FA_X1 U1294 ( .A(n1854), .B(n1873), .CI(n1856), .CO(n1849), .S(n1850) );
  FA_X1 U1295 ( .A(n1877), .B(n1879), .CI(n1875), .CO(n1851), .S(n1852) );
  FA_X1 U1296 ( .A(n2455), .B(n2519), .CI(n2487), .CO(n1853), .S(n1854) );
  FA_X1 U1297 ( .A(n2391), .B(n2551), .CI(n2423), .CO(n1855), .S(n1856) );
  FA_X1 U1298 ( .A(n2327), .B(n2583), .CI(n2359), .CO(n1857), .S(n1858) );
  FA_X1 U1299 ( .A(n2295), .B(n2615), .CI(n2263), .CO(n1859), .S(n1860) );
  FA_X1 U1300 ( .A(n1883), .B(n1866), .CI(n1864), .CO(n1861), .S(n1862) );
  FA_X1 U1301 ( .A(n1868), .B(n1870), .CI(n1885), .CO(n1863), .S(n1864) );
  FA_X1 U1302 ( .A(n1872), .B(n1889), .CI(n1887), .CO(n1865), .S(n1866) );
  FA_X1 U1303 ( .A(n1878), .B(n1874), .CI(n1876), .CO(n1867), .S(n1868) );
  FA_X1 U1304 ( .A(n1893), .B(n1895), .CI(n1891), .CO(n1869), .S(n1870) );
  FA_X1 U1305 ( .A(n1880), .B(n2488), .CI(n1897), .CO(n1871), .S(n1872) );
  FA_X1 U1306 ( .A(n2360), .B(n2520), .CI(n2392), .CO(n1873), .S(n1874) );
  FA_X1 U1307 ( .A(n2328), .B(n2552), .CI(n2424), .CO(n1875), .S(n1876) );
  FA_X1 U1308 ( .A(n2616), .B(n2456), .CI(n2584), .CO(n1877), .S(n1878) );
  HA_X1 U1309 ( .A(n2296), .B(n2066), .CO(n1879), .S(n1880) );
  FA_X1 U1310 ( .A(n1901), .B(n1886), .CI(n1884), .CO(n1881), .S(n1882) );
  FA_X1 U1311 ( .A(n1888), .B(n1890), .CI(n1903), .CO(n1883), .S(n1884) );
  FA_X1 U1312 ( .A(n1907), .B(n1892), .CI(n1905), .CO(n1885), .S(n1886) );
  FA_X1 U1313 ( .A(n1898), .B(n1894), .CI(n1896), .CO(n1887), .S(n1888) );
  FA_X1 U1314 ( .A(n1909), .B(n1913), .CI(n1911), .CO(n1889), .S(n1890) );
  FA_X1 U1315 ( .A(n2489), .B(n2521), .CI(n1915), .CO(n1891), .S(n1892) );
  FA_X1 U1316 ( .A(n2425), .B(n2553), .CI(n2457), .CO(n1893), .S(n1894) );
  FA_X1 U1317 ( .A(n2361), .B(n2585), .CI(n2393), .CO(n1895), .S(n1896) );
  FA_X1 U1318 ( .A(n2297), .B(n2617), .CI(n2329), .CO(n1897), .S(n1898) );
  FA_X1 U1319 ( .A(n1919), .B(n1904), .CI(n1902), .CO(n1899), .S(n1900) );
  FA_X1 U1320 ( .A(n1906), .B(n1923), .CI(n1921), .CO(n1901), .S(n1902) );
  FA_X1 U1321 ( .A(n1925), .B(n1914), .CI(n1908), .CO(n1903), .S(n1904) );
  FA_X1 U1322 ( .A(n1910), .B(n1927), .CI(n1912), .CO(n1905), .S(n1906) );
  FA_X1 U1323 ( .A(n1931), .B(n1916), .CI(n1929), .CO(n1907), .S(n1908) );
  FA_X1 U1324 ( .A(n2458), .B(n2586), .CI(n2554), .CO(n1909), .S(n1910) );
  FA_X1 U1325 ( .A(n2618), .B(n2522), .CI(n2426), .CO(n1911), .S(n1912) );
  FA_X1 U1326 ( .A(n2362), .B(n2490), .CI(n2394), .CO(n1913), .S(n1914) );
  HA_X1 U1327 ( .A(n2330), .B(n2067), .CO(n1915), .S(n1916) );
  FA_X1 U1328 ( .A(n1935), .B(n1922), .CI(n1920), .CO(n1917), .S(n1918) );
  FA_X1 U1329 ( .A(n1924), .B(n1926), .CI(n1937), .CO(n1919), .S(n1920) );
  FA_X1 U1330 ( .A(n1941), .B(n1932), .CI(n1939), .CO(n1921), .S(n1922) );
  FA_X1 U1331 ( .A(n1928), .B(n1943), .CI(n1930), .CO(n1923), .S(n1924) );
  FA_X1 U1332 ( .A(n1947), .B(n2523), .CI(n1945), .CO(n1925), .S(n1926) );
  FA_X1 U1333 ( .A(n2459), .B(n2555), .CI(n2491), .CO(n1927), .S(n1928) );
  FA_X1 U1334 ( .A(n2395), .B(n2587), .CI(n2427), .CO(n1929), .S(n1930) );
  FA_X1 U1335 ( .A(n2363), .B(n2619), .CI(n2331), .CO(n1931), .S(n1932) );
  FA_X1 U1336 ( .A(n1938), .B(n1951), .CI(n1936), .CO(n1933), .S(n1934) );
  FA_X1 U1337 ( .A(n1953), .B(n1942), .CI(n1940), .CO(n1935), .S(n1936) );
  FA_X1 U1338 ( .A(n1946), .B(n1944), .CI(n1955), .CO(n1937), .S(n1938) );
  FA_X1 U1339 ( .A(n1957), .B(n1961), .CI(n1959), .CO(n1939), .S(n1940) );
  FA_X1 U1340 ( .A(n2556), .B(n2588), .CI(n1948), .CO(n1941), .S(n1942) );
  FA_X1 U1341 ( .A(n2428), .B(n2524), .CI(n2460), .CO(n1943), .S(n1944) );
  FA_X1 U1342 ( .A(n2396), .B(n2492), .CI(n2620), .CO(n1945), .S(n1946) );
  HA_X1 U1343 ( .A(n2364), .B(n2068), .CO(n1947), .S(n1948) );
  FA_X1 U1344 ( .A(n1965), .B(n1954), .CI(n1952), .CO(n1949), .S(n1950) );
  FA_X1 U1345 ( .A(n1967), .B(n1969), .CI(n1956), .CO(n1951), .S(n1952) );
  FA_X1 U1346 ( .A(n1960), .B(n1962), .CI(n1958), .CO(n1953), .S(n1954) );
  FA_X1 U1347 ( .A(n1973), .B(n1975), .CI(n1971), .CO(n1955), .S(n1956) );
  FA_X1 U1348 ( .A(n2493), .B(n2557), .CI(n2525), .CO(n1957), .S(n1958) );
  FA_X1 U1349 ( .A(n2429), .B(n2589), .CI(n2461), .CO(n1959), .S(n1960) );
  FA_X1 U1350 ( .A(n2397), .B(n2621), .CI(n2365), .CO(n1961), .S(n1962) );
  FA_X1 U1351 ( .A(n1979), .B(n1968), .CI(n1966), .CO(n1963), .S(n1964) );
  FA_X1 U1352 ( .A(n1981), .B(n1974), .CI(n1970), .CO(n1965), .S(n1966) );
  FA_X1 U1353 ( .A(n1983), .B(n1985), .CI(n1972), .CO(n1967), .S(n1968) );
  FA_X1 U1354 ( .A(n1976), .B(n2494), .CI(n1987), .CO(n1969), .S(n1970) );
  FA_X1 U1355 ( .A(n2558), .B(n2430), .CI(n2462), .CO(n1971), .S(n1972) );
  FA_X1 U1356 ( .A(n2622), .B(n2526), .CI(n2590), .CO(n1973), .S(n1974) );
  HA_X1 U1357 ( .A(n2398), .B(n2069), .CO(n1975), .S(n1976) );
  FA_X1 U1358 ( .A(n1991), .B(n1982), .CI(n1980), .CO(n1977), .S(n1978) );
  FA_X1 U1359 ( .A(n1984), .B(n1988), .CI(n1993), .CO(n1979), .S(n1980) );
  FA_X1 U1360 ( .A(n1995), .B(n1997), .CI(n1986), .CO(n1981), .S(n1982) );
  FA_X1 U1361 ( .A(n2527), .B(n2559), .CI(n1999), .CO(n1983), .S(n1984) );
  FA_X1 U1362 ( .A(n2463), .B(n2591), .CI(n2495), .CO(n1985), .S(n1986) );
  FA_X1 U1363 ( .A(n2431), .B(n2623), .CI(n2399), .CO(n1987), .S(n1988) );
  FA_X1 U1364 ( .A(n2003), .B(n1994), .CI(n1992), .CO(n1989), .S(n1990) );
  FA_X1 U1365 ( .A(n1998), .B(n1996), .CI(n2005), .CO(n1991), .S(n1992) );
  FA_X1 U1366 ( .A(n2009), .B(n2000), .CI(n2007), .CO(n1993), .S(n1994) );
  FA_X1 U1367 ( .A(n2464), .B(n2560), .CI(n2496), .CO(n1995), .S(n1996) );
  FA_X1 U1368 ( .A(n2624), .B(n2528), .CI(n2592), .CO(n1997), .S(n1998) );
  HA_X1 U1369 ( .A(n2432), .B(n2070), .CO(n1999), .S(n2000) );
  FA_X1 U1370 ( .A(n2006), .B(n2013), .CI(n2004), .CO(n2001), .S(n2002) );
  FA_X1 U1371 ( .A(n2010), .B(n2008), .CI(n2015), .CO(n2003), .S(n2004) );
  FA_X1 U1372 ( .A(n2019), .B(n2561), .CI(n2017), .CO(n2005), .S(n2006) );
  FA_X1 U1373 ( .A(n2497), .B(n2593), .CI(n2529), .CO(n2007), .S(n2008) );
  FA_X1 U1374 ( .A(n2465), .B(n2625), .CI(n2433), .CO(n2009), .S(n2010) );
  FA_X1 U1375 ( .A(n2023), .B(n2016), .CI(n2014), .CO(n2011), .S(n2012) );
  FA_X1 U1376 ( .A(n2025), .B(n2027), .CI(n2018), .CO(n2013), .S(n2014) );
  FA_X1 U1377 ( .A(n2498), .B(n2530), .CI(n2020), .CO(n2015), .S(n2016) );
  FA_X1 U1378 ( .A(n2626), .B(n2562), .CI(n2594), .CO(n2017), .S(n2018) );
  HA_X1 U1379 ( .A(n2466), .B(n2071), .CO(n2019), .S(n2020) );
  FA_X1 U1380 ( .A(n2031), .B(n2028), .CI(n2024), .CO(n2021), .S(n2022) );
  FA_X1 U1381 ( .A(n2033), .B(n2035), .CI(n2026), .CO(n2023), .S(n2024) );
  FA_X1 U1382 ( .A(n2531), .B(n2595), .CI(n2563), .CO(n2025), .S(n2026) );
  FA_X1 U1383 ( .A(n2499), .B(n2627), .CI(n2467), .CO(n2027), .S(n2028) );
  FA_X1 U1384 ( .A(n2034), .B(n2039), .CI(n2032), .CO(n2029), .S(n2030) );
  FA_X1 U1385 ( .A(n2036), .B(n2628), .CI(n2041), .CO(n2031), .S(n2032) );
  FA_X1 U1386 ( .A(n2532), .B(n2564), .CI(n2596), .CO(n2033), .S(n2034) );
  HA_X1 U1387 ( .A(n2500), .B(n2072), .CO(n2035), .S(n2036) );
  FA_X1 U1388 ( .A(n2042), .B(n2045), .CI(n2040), .CO(n2037), .S(n2038) );
  FA_X1 U1389 ( .A(n2565), .B(n2597), .CI(n2047), .CO(n2039), .S(n2040) );
  FA_X1 U1390 ( .A(n2533), .B(n2629), .CI(n2501), .CO(n2041), .S(n2042) );
  FA_X1 U1391 ( .A(n2051), .B(n2048), .CI(n2046), .CO(n2043), .S(n2044) );
  FA_X1 U1392 ( .A(n2566), .B(n2630), .CI(n2598), .CO(n2045), .S(n2046) );
  HA_X1 U1393 ( .A(n2534), .B(n2073), .CO(n2047), .S(n2048) );
  FA_X1 U1394 ( .A(n2055), .B(n2599), .CI(n2052), .CO(n2049), .S(n2050) );
  FA_X1 U1395 ( .A(n2567), .B(n2631), .CI(n2535), .CO(n2051), .S(n2052) );
  FA_X1 U1396 ( .A(n2600), .B(n2632), .CI(n2056), .CO(n2053), .S(n2054) );
  HA_X1 U1397 ( .A(n2568), .B(n2074), .CO(n2055), .S(n2056) );
  FA_X1 U1398 ( .A(n2601), .B(n2633), .CI(n2569), .CO(n2057), .S(n2058) );
  HA_X1 U1399 ( .A(n2634), .B(n2602), .CO(n2059), .S(n2060) );
  NOR2_X4 U1400 ( .A1(n2637), .A2(n3575), .ZN(n2077) );
  NOR2_X4 U1401 ( .A1(n2638), .A2(n3575), .ZN(n1044) );
  NOR2_X4 U1402 ( .A1(n2639), .A2(n3575), .ZN(n2078) );
  NOR2_X4 U1403 ( .A1(n2640), .A2(n3575), .ZN(n1054) );
  NOR2_X4 U1404 ( .A1(n2641), .A2(n3575), .ZN(n2079) );
  NOR2_X4 U1405 ( .A1(n2642), .A2(n3575), .ZN(n1068) );
  NOR2_X4 U1406 ( .A1(n2643), .A2(n3575), .ZN(n2080) );
  NOR2_X4 U1407 ( .A1(n2644), .A2(n3575), .ZN(n1086) );
  NOR2_X4 U1408 ( .A1(n2645), .A2(n3575), .ZN(n2081) );
  NOR2_X4 U1409 ( .A1(n2646), .A2(n3575), .ZN(n1108) );
  NOR2_X4 U1410 ( .A1(n2647), .A2(n3575), .ZN(n2082) );
  NOR2_X4 U1411 ( .A1(n2648), .A2(n3575), .ZN(n1134) );
  NOR2_X4 U1412 ( .A1(n2649), .A2(n3575), .ZN(n2083) );
  NOR2_X4 U1413 ( .A1(n2650), .A2(n3575), .ZN(n1164) );
  NOR2_X4 U1414 ( .A1(n2651), .A2(n3575), .ZN(n2084) );
  NOR2_X4 U1415 ( .A1(n2652), .A2(n3575), .ZN(n1198) );
  NOR2_X4 U1416 ( .A1(n2653), .A2(n3575), .ZN(n2085) );
  NOR2_X4 U1417 ( .A1(n2654), .A2(n3575), .ZN(n1236) );
  NOR2_X4 U1418 ( .A1(n2655), .A2(n3575), .ZN(n2086) );
  NOR2_X4 U1419 ( .A1(n2656), .A2(n3575), .ZN(n1278) );
  NOR2_X4 U1420 ( .A1(n2657), .A2(n3575), .ZN(n2087) );
  NOR2_X4 U1421 ( .A1(n2658), .A2(n3575), .ZN(n1324) );
  NOR2_X4 U1422 ( .A1(n2659), .A2(n3575), .ZN(n2088) );
  NOR2_X4 U1423 ( .A1(n2660), .A2(n3575), .ZN(n1374) );
  NOR2_X4 U1424 ( .A1(n2661), .A2(n3575), .ZN(n2089) );
  NOR2_X4 U1425 ( .A1(n2662), .A2(n3575), .ZN(n1428) );
  NOR2_X4 U1426 ( .A1(n2663), .A2(n3575), .ZN(n2090) );
  NOR2_X4 U1427 ( .A1(n2664), .A2(n3575), .ZN(n1486) );
  NOR2_X4 U1428 ( .A1(n2665), .A2(n3575), .ZN(n2091) );
  NOR2_X4 U1429 ( .A1(n2666), .A2(n3575), .ZN(n2092) );
  NOR2_X4 U1430 ( .A1(n2667), .A2(n3575), .ZN(n1548) );
  OAI22_X2 U1463 ( .A1(n3458), .A2(n2668), .B1(n3642), .B2(n3575), .ZN(n2095)
         );
  OAI22_X2 U1464 ( .A1(n3458), .A2(n2669), .B1(n2668), .B2(n3642), .ZN(n2096)
         );
  OAI22_X2 U1465 ( .A1(n3458), .A2(n2670), .B1(n2669), .B2(n3642), .ZN(n2097)
         );
  OAI22_X2 U1466 ( .A1(n3458), .A2(n2671), .B1(n2670), .B2(n3642), .ZN(n2098)
         );
  OAI22_X2 U1467 ( .A1(n3458), .A2(n2672), .B1(n2671), .B2(n3642), .ZN(n2099)
         );
  OAI22_X2 U1468 ( .A1(n3458), .A2(n2673), .B1(n2672), .B2(n3642), .ZN(n2100)
         );
  OAI22_X2 U1469 ( .A1(n3458), .A2(n2674), .B1(n2673), .B2(n3642), .ZN(n2101)
         );
  OAI22_X2 U1470 ( .A1(n3458), .A2(n2675), .B1(n2674), .B2(n3642), .ZN(n2102)
         );
  OAI22_X2 U1471 ( .A1(n3458), .A2(n2676), .B1(n2675), .B2(n3642), .ZN(n2103)
         );
  OAI22_X2 U1472 ( .A1(n3458), .A2(n2677), .B1(n2676), .B2(n3642), .ZN(n2104)
         );
  OAI22_X2 U1473 ( .A1(n3458), .A2(n2678), .B1(n2677), .B2(n3642), .ZN(n2105)
         );
  OAI22_X2 U1474 ( .A1(n3458), .A2(n2679), .B1(n2678), .B2(n3642), .ZN(n2106)
         );
  OAI22_X2 U1475 ( .A1(n3458), .A2(n2680), .B1(n2679), .B2(n3642), .ZN(n2107)
         );
  OAI22_X2 U1476 ( .A1(n3458), .A2(n2681), .B1(n2680), .B2(n3642), .ZN(n2108)
         );
  OAI22_X2 U1478 ( .A1(n3458), .A2(n2683), .B1(n2682), .B2(n3642), .ZN(n2110)
         );
  OAI22_X2 U1479 ( .A1(n3458), .A2(n2684), .B1(n2683), .B2(n3642), .ZN(n2111)
         );
  OAI22_X2 U1480 ( .A1(n3458), .A2(n2685), .B1(n2684), .B2(n3642), .ZN(n2112)
         );
  OAI22_X2 U1481 ( .A1(n3458), .A2(n2686), .B1(n2685), .B2(n3642), .ZN(n2113)
         );
  OAI22_X2 U1482 ( .A1(n3457), .A2(n2687), .B1(n2686), .B2(n3642), .ZN(n2114)
         );
  OAI22_X2 U1483 ( .A1(n3458), .A2(n2688), .B1(n2687), .B2(n3642), .ZN(n2115)
         );
  OAI22_X2 U1484 ( .A1(n3458), .A2(n2689), .B1(n2688), .B2(n3642), .ZN(n2116)
         );
  OAI22_X2 U1485 ( .A1(n3458), .A2(n2690), .B1(n2689), .B2(n3642), .ZN(n2117)
         );
  OAI22_X2 U1487 ( .A1(n3458), .A2(n2692), .B1(n2691), .B2(n3642), .ZN(n2119)
         );
  OAI22_X2 U1594 ( .A1(n3614), .A2(n2735), .B1(n2734), .B2(n3742), .ZN(n2164)
         );
  OAI22_X2 U1595 ( .A1(n3614), .A2(n2736), .B1(n2735), .B2(n3742), .ZN(n2165)
         );
  OAI22_X2 U1596 ( .A1(n3614), .A2(n2737), .B1(n2736), .B2(n3741), .ZN(n2166)
         );
  OAI22_X2 U1597 ( .A1(n3614), .A2(n2738), .B1(n2737), .B2(n3742), .ZN(n2167)
         );
  OAI22_X2 U1598 ( .A1(n3614), .A2(n2739), .B1(n2738), .B2(n3741), .ZN(n2168)
         );
  OAI22_X2 U1599 ( .A1(n3614), .A2(n2740), .B1(n2739), .B2(n3742), .ZN(n2169)
         );
  OAI22_X2 U1600 ( .A1(n3614), .A2(n2741), .B1(n2740), .B2(n3741), .ZN(n2170)
         );
  OAI22_X2 U1601 ( .A1(n3614), .A2(n2742), .B1(n2741), .B2(n3741), .ZN(n2171)
         );
  OAI22_X2 U1602 ( .A1(n3614), .A2(n2743), .B1(n2742), .B2(n3741), .ZN(n2172)
         );
  OAI22_X2 U1603 ( .A1(n3614), .A2(n2744), .B1(n2743), .B2(n3742), .ZN(n2173)
         );
  OAI22_X2 U1604 ( .A1(n3614), .A2(n2745), .B1(n2744), .B2(n3741), .ZN(n2174)
         );
  OAI22_X2 U1606 ( .A1(n3614), .A2(n2747), .B1(n2746), .B2(n3742), .ZN(n2176)
         );
  OAI22_X2 U1608 ( .A1(n3614), .A2(n2749), .B1(n2748), .B2(n3742), .ZN(n2178)
         );
  OAI22_X2 U1609 ( .A1(n3614), .A2(n2750), .B1(n2749), .B2(n3741), .ZN(n2179)
         );
  OAI22_X2 U1610 ( .A1(n3614), .A2(n2751), .B1(n2750), .B2(n3742), .ZN(n2180)
         );
  OAI22_X2 U1611 ( .A1(n3614), .A2(n2752), .B1(n2751), .B2(n3741), .ZN(n2181)
         );
  OAI22_X2 U1658 ( .A1(n3706), .A2(n2767), .B1(n3581), .B2(n3280), .ZN(n2197)
         );
  OAI22_X2 U1659 ( .A1(n3705), .A2(n2768), .B1(n2767), .B2(n3581), .ZN(n2198)
         );
  OAI22_X2 U1660 ( .A1(n3706), .A2(n2769), .B1(n2768), .B2(n3581), .ZN(n2199)
         );
  OAI22_X2 U1661 ( .A1(n3706), .A2(n2770), .B1(n2769), .B2(n3581), .ZN(n2200)
         );
  OAI22_X2 U1662 ( .A1(n3705), .A2(n2771), .B1(n2770), .B2(n3581), .ZN(n2201)
         );
  OAI22_X2 U1663 ( .A1(n3705), .A2(n2772), .B1(n2771), .B2(n3581), .ZN(n2202)
         );
  OAI22_X2 U1664 ( .A1(n3705), .A2(n2773), .B1(n2772), .B2(n3581), .ZN(n2203)
         );
  OAI22_X2 U1665 ( .A1(n3706), .A2(n2774), .B1(n2773), .B2(n3581), .ZN(n2204)
         );
  OAI22_X2 U1666 ( .A1(n3705), .A2(n2775), .B1(n2774), .B2(n3581), .ZN(n2205)
         );
  OAI22_X2 U1667 ( .A1(n3705), .A2(n2776), .B1(n2775), .B2(n3581), .ZN(n2206)
         );
  OAI22_X2 U1668 ( .A1(n3705), .A2(n2777), .B1(n2776), .B2(n3581), .ZN(n2207)
         );
  OAI22_X2 U1669 ( .A1(n3706), .A2(n2778), .B1(n2777), .B2(n3581), .ZN(n2208)
         );
  OAI22_X2 U1670 ( .A1(n3706), .A2(n2779), .B1(n2778), .B2(n3581), .ZN(n2209)
         );
  OAI22_X2 U1671 ( .A1(n3705), .A2(n2780), .B1(n2779), .B2(n3581), .ZN(n2210)
         );
  OAI22_X2 U1672 ( .A1(n3706), .A2(n2781), .B1(n2780), .B2(n3581), .ZN(n2211)
         );
  OAI22_X2 U1673 ( .A1(n3705), .A2(n2782), .B1(n2781), .B2(n3581), .ZN(n2212)
         );
  OAI22_X2 U1674 ( .A1(n3705), .A2(n2783), .B1(n2782), .B2(n3581), .ZN(n2213)
         );
  OAI22_X2 U1677 ( .A1(n3705), .A2(n2786), .B1(n2785), .B2(n3581), .ZN(n2216)
         );
  OAI22_X2 U1678 ( .A1(n3705), .A2(n2787), .B1(n2786), .B2(n3581), .ZN(n2217)
         );
  OAI22_X2 U1682 ( .A1(n3705), .A2(n2791), .B1(n2790), .B2(n3581), .ZN(n2221)
         );
  OAI22_X2 U1683 ( .A1(n3705), .A2(n2792), .B1(n2791), .B2(n3581), .ZN(n2222)
         );
  OAI22_X2 U1685 ( .A1(n3706), .A2(n2794), .B1(n3581), .B2(n2793), .ZN(n2224)
         );
  OAI22_X2 U1686 ( .A1(n3705), .A2(n2795), .B1(n2794), .B2(n3581), .ZN(n2225)
         );
  OAI22_X2 U1687 ( .A1(n3706), .A2(n2796), .B1(n2795), .B2(n3581), .ZN(n2226)
         );
  OAI22_X2 U1688 ( .A1(n3706), .A2(n2797), .B1(n2796), .B2(n3581), .ZN(n2227)
         );
  OAI22_X2 U1854 ( .A1(n3491), .A2(n2867), .B1(n2866), .B2(n3729), .ZN(n2300)
         );
  OAI22_X2 U1855 ( .A1(n3491), .A2(n2868), .B1(n2867), .B2(n3729), .ZN(n2301)
         );
  OAI22_X2 U1856 ( .A1(n3491), .A2(n2869), .B1(n2868), .B2(n3729), .ZN(n2302)
         );
  OAI22_X2 U1857 ( .A1(n3491), .A2(n2870), .B1(n2869), .B2(n3729), .ZN(n2303)
         );
  OAI22_X2 U1858 ( .A1(n3491), .A2(n2871), .B1(n2870), .B2(n3728), .ZN(n2304)
         );
  OAI22_X2 U1859 ( .A1(n3491), .A2(n2872), .B1(n2871), .B2(n3728), .ZN(n2305)
         );
  OAI22_X2 U1860 ( .A1(n3491), .A2(n2873), .B1(n2872), .B2(n3729), .ZN(n2306)
         );
  OAI22_X2 U1861 ( .A1(n3491), .A2(n2874), .B1(n2873), .B2(n3728), .ZN(n2307)
         );
  OAI22_X2 U1862 ( .A1(n3491), .A2(n2875), .B1(n2874), .B2(n3728), .ZN(n2308)
         );
  OAI22_X2 U1863 ( .A1(n3491), .A2(n2876), .B1(n2875), .B2(n3729), .ZN(n2309)
         );
  OAI22_X2 U1865 ( .A1(n3491), .A2(n2878), .B1(n2877), .B2(n3728), .ZN(n2311)
         );
  OAI22_X2 U1872 ( .A1(n3491), .A2(n2885), .B1(n2884), .B2(n3728), .ZN(n2318)
         );
  OAI22_X2 U1873 ( .A1(n3491), .A2(n2886), .B1(n2885), .B2(n3729), .ZN(n2319)
         );
  OAI22_X2 U1874 ( .A1(n3491), .A2(n2887), .B1(n2886), .B2(n3729), .ZN(n2320)
         );
  OAI22_X2 U1876 ( .A1(n3491), .A2(n2889), .B1(n2888), .B2(n3728), .ZN(n2322)
         );
  OAI22_X2 U1878 ( .A1(n3491), .A2(n2891), .B1(n2890), .B2(n3728), .ZN(n2324)
         );
  OAI22_X2 U1880 ( .A1(n3491), .A2(n2893), .B1(n2892), .B2(n3728), .ZN(n2326)
         );
  OAI22_X2 U1881 ( .A1(n3491), .A2(n2894), .B1(n2893), .B2(n3729), .ZN(n2327)
         );
  OAI22_X2 U1927 ( .A1(n443), .A2(n2908), .B1(n2907), .B2(n393), .ZN(n2342) );
  OAI22_X2 U1932 ( .A1(n443), .A2(n2913), .B1(n2912), .B2(n393), .ZN(n2347) );
  OAI22_X2 U1982 ( .A1(n3578), .A2(n3285), .B1(n2964), .B2(n3625), .ZN(n2069)
         );
  OAI22_X2 U1983 ( .A1(n3578), .A2(n2932), .B1(n3625), .B2(n3285), .ZN(n2367)
         );
  OAI22_X2 U1984 ( .A1(n3578), .A2(n2933), .B1(n2932), .B2(n3626), .ZN(n2368)
         );
  OAI22_X2 U1985 ( .A1(n3578), .A2(n2934), .B1(n2933), .B2(n3626), .ZN(n2369)
         );
  OAI22_X2 U1986 ( .A1(n3578), .A2(n2935), .B1(n2934), .B2(n3626), .ZN(n2370)
         );
  OAI22_X2 U1987 ( .A1(n3578), .A2(n2936), .B1(n2935), .B2(n3625), .ZN(n2371)
         );
  OAI22_X2 U1988 ( .A1(n3578), .A2(n2937), .B1(n2936), .B2(n3625), .ZN(n2372)
         );
  OAI22_X2 U1989 ( .A1(n3578), .A2(n2938), .B1(n2937), .B2(n3626), .ZN(n2373)
         );
  OAI22_X2 U1990 ( .A1(n440), .A2(n2939), .B1(n2938), .B2(n3626), .ZN(n2374)
         );
  OAI22_X2 U1991 ( .A1(n3578), .A2(n2940), .B1(n2939), .B2(n3626), .ZN(n2375)
         );
  OAI22_X2 U1992 ( .A1(n3578), .A2(n2941), .B1(n2940), .B2(n3625), .ZN(n2376)
         );
  OAI22_X2 U1993 ( .A1(n440), .A2(n2942), .B1(n2941), .B2(n3625), .ZN(n2377)
         );
  OAI22_X2 U1994 ( .A1(n440), .A2(n2943), .B1(n2942), .B2(n3625), .ZN(n2378)
         );
  OAI22_X2 U1995 ( .A1(n3578), .A2(n2944), .B1(n2943), .B2(n3625), .ZN(n2379)
         );
  OAI22_X2 U1996 ( .A1(n440), .A2(n2945), .B1(n2944), .B2(n3626), .ZN(n2380)
         );
  OAI22_X2 U1997 ( .A1(n3578), .A2(n2946), .B1(n2945), .B2(n3626), .ZN(n2381)
         );
  OAI22_X2 U1998 ( .A1(n3578), .A2(n2947), .B1(n2946), .B2(n3626), .ZN(n2382)
         );
  OAI22_X2 U1999 ( .A1(n440), .A2(n2948), .B1(n2947), .B2(n3626), .ZN(n2383)
         );
  OAI22_X2 U2001 ( .A1(n440), .A2(n2950), .B1(n2949), .B2(n3625), .ZN(n2385)
         );
  OAI22_X2 U2002 ( .A1(n440), .A2(n2951), .B1(n2950), .B2(n3625), .ZN(n2386)
         );
  OAI22_X2 U2003 ( .A1(n440), .A2(n2952), .B1(n2951), .B2(n3625), .ZN(n2387)
         );
  OAI22_X2 U2004 ( .A1(n3578), .A2(n2953), .B1(n2952), .B2(n3626), .ZN(n2388)
         );
  OAI22_X2 U2005 ( .A1(n440), .A2(n2954), .B1(n2953), .B2(n3626), .ZN(n2389)
         );
  OAI22_X2 U2006 ( .A1(n3578), .A2(n2955), .B1(n2954), .B2(n3625), .ZN(n2390)
         );
  OAI22_X2 U2007 ( .A1(n3578), .A2(n2956), .B1(n2955), .B2(n3625), .ZN(n2391)
         );
  OAI22_X2 U2008 ( .A1(n3578), .A2(n2957), .B1(n2956), .B2(n3625), .ZN(n2392)
         );
  OAI22_X2 U2009 ( .A1(n3578), .A2(n2958), .B1(n2957), .B2(n3625), .ZN(n2393)
         );
  OAI22_X2 U2010 ( .A1(n3578), .A2(n2959), .B1(n2958), .B2(n3626), .ZN(n2394)
         );
  OAI22_X2 U2011 ( .A1(n440), .A2(n2960), .B1(n2959), .B2(n3626), .ZN(n2395)
         );
  OAI22_X2 U2012 ( .A1(n3578), .A2(n2961), .B1(n2960), .B2(n3625), .ZN(n2396)
         );
  OAI22_X2 U2013 ( .A1(n440), .A2(n2962), .B1(n2961), .B2(n3626), .ZN(n2397)
         );
  OAI22_X2 U2014 ( .A1(n3578), .A2(n2963), .B1(n2962), .B2(n3626), .ZN(n2398)
         );
  OAI22_X2 U2251 ( .A1(n3620), .A2(n3072), .B1(n3071), .B2(n3679), .ZN(n2511)
         );
  OAI22_X2 U2258 ( .A1(n3620), .A2(n3079), .B1(n3078), .B2(n3679), .ZN(n2518)
         );
  OAI22_X2 U2259 ( .A1(n428), .A2(n3080), .B1(n3079), .B2(n3679), .ZN(n2519)
         );
  OAI22_X2 U2267 ( .A1(n3620), .A2(n3088), .B1(n3087), .B2(n3679), .ZN(n2527)
         );
  OAI22_X2 U2272 ( .A1(n3620), .A2(n3093), .B1(n3092), .B2(n3679), .ZN(n2532)
         );
  OAI22_X2 U2273 ( .A1(n3620), .A2(n3094), .B1(n3093), .B2(n3679), .ZN(n2533)
         );
  OAI22_X2 U2307 ( .A1(n3712), .A2(n3290), .B1(n3129), .B2(n3674), .ZN(n2074)
         );
  OAI22_X2 U2312 ( .A1(n425), .A2(n3101), .B1(n3100), .B2(n3674), .ZN(n2541)
         );
  OAI22_X2 U2316 ( .A1(n425), .A2(n3105), .B1(n3104), .B2(n3674), .ZN(n2545)
         );
  OAI22_X2 U2317 ( .A1(n425), .A2(n3106), .B1(n3105), .B2(n3674), .ZN(n2546)
         );
  OAI22_X2 U2319 ( .A1(n425), .A2(n3108), .B1(n3107), .B2(n3674), .ZN(n2548)
         );
  OAI22_X2 U2320 ( .A1(n425), .A2(n3109), .B1(n3108), .B2(n3674), .ZN(n2549)
         );
  OAI22_X2 U2321 ( .A1(n425), .A2(n3110), .B1(n3109), .B2(n3674), .ZN(n2550)
         );
  OAI22_X2 U2323 ( .A1(n425), .A2(n3112), .B1(n3111), .B2(n3674), .ZN(n2552)
         );
  OAI22_X2 U2327 ( .A1(n3712), .A2(n3116), .B1(n3115), .B2(n3674), .ZN(n2556)
         );
  OAI22_X2 U2328 ( .A1(n425), .A2(n3117), .B1(n3116), .B2(n3674), .ZN(n2557)
         );
  OAI22_X2 U2330 ( .A1(n425), .A2(n3119), .B1(n3118), .B2(n3674), .ZN(n2559)
         );
  OAI22_X2 U2331 ( .A1(n425), .A2(n3120), .B1(n3119), .B2(n3674), .ZN(n2560)
         );
  OAI22_X2 U2332 ( .A1(n3712), .A2(n3121), .B1(n3120), .B2(n3674), .ZN(n2561)
         );
  OAI22_X2 U2333 ( .A1(n425), .A2(n3122), .B1(n3121), .B2(n3674), .ZN(n2562)
         );
  OAI22_X2 U2334 ( .A1(n3712), .A2(n3123), .B1(n3122), .B2(n3674), .ZN(n2563)
         );
  OAI22_X2 U2335 ( .A1(n3712), .A2(n3124), .B1(n3123), .B2(n3674), .ZN(n2564)
         );
  OAI22_X2 U2336 ( .A1(n3712), .A2(n3125), .B1(n3124), .B2(n3674), .ZN(n2565)
         );
  OAI22_X2 U2337 ( .A1(n3712), .A2(n3126), .B1(n3125), .B2(n3674), .ZN(n2566)
         );
  OAI22_X2 U2339 ( .A1(n3712), .A2(n3128), .B1(n3127), .B2(n3674), .ZN(n2568)
         );
  OAI22_X2 U2375 ( .A1(n3722), .A2(n3132), .B1(n3131), .B2(n3573), .ZN(n2573)
         );
  OAI22_X2 U2377 ( .A1(n3722), .A2(n3134), .B1(n3133), .B2(n372), .ZN(n2575)
         );
  OAI22_X2 U2380 ( .A1(n3722), .A2(n3137), .B1(n3136), .B2(n3573), .ZN(n2578)
         );
  OAI22_X2 U2385 ( .A1(n3722), .A2(n3142), .B1(n3141), .B2(n3573), .ZN(n2583)
         );
  OAI22_X2 U2386 ( .A1(n3722), .A2(n3143), .B1(n3142), .B2(n3573), .ZN(n2584)
         );
  OAI22_X2 U2388 ( .A1(n3722), .A2(n3145), .B1(n3144), .B2(n372), .ZN(n2586)
         );
  OAI22_X2 U2389 ( .A1(n3722), .A2(n3146), .B1(n3145), .B2(n3573), .ZN(n2587)
         );
  OAI22_X2 U2396 ( .A1(n3722), .A2(n3153), .B1(n3152), .B2(n3573), .ZN(n2594)
         );
  OAI22_X2 U2399 ( .A1(n3722), .A2(n3156), .B1(n3155), .B2(n3573), .ZN(n2597)
         );
  OAI22_X2 U2402 ( .A1(n3722), .A2(n3159), .B1(n3158), .B2(n3573), .ZN(n2600)
         );
  OAI22_X2 U2404 ( .A1(n3722), .A2(n3161), .B1(n3160), .B2(n3573), .ZN(n2602)
         );
  OAI22_X2 U2441 ( .A1(n419), .A2(n3166), .B1(n3165), .B2(n369), .ZN(n2608) );
  OAI22_X2 U2442 ( .A1(n419), .A2(n3167), .B1(n3166), .B2(n369), .ZN(n2609) );
  OAI22_X2 U2444 ( .A1(n419), .A2(n3169), .B1(n3168), .B2(n369), .ZN(n2611) );
  OAI22_X2 U2445 ( .A1(n419), .A2(n3170), .B1(n3169), .B2(n369), .ZN(n2612) );
  OAI22_X2 U2446 ( .A1(n419), .A2(n3171), .B1(n3170), .B2(n369), .ZN(n2613) );
  OAI22_X2 U2447 ( .A1(n419), .A2(n3172), .B1(n3171), .B2(n369), .ZN(n2614) );
  OAI22_X2 U2448 ( .A1(n419), .A2(n3173), .B1(n3172), .B2(n369), .ZN(n2615) );
  OAI22_X2 U2449 ( .A1(n419), .A2(n3174), .B1(n3173), .B2(n369), .ZN(n2616) );
  OAI22_X2 U2450 ( .A1(n419), .A2(n3175), .B1(n3174), .B2(n369), .ZN(n2617) );
  OAI22_X2 U2452 ( .A1(n419), .A2(n3177), .B1(n3176), .B2(n369), .ZN(n2619) );
  OAI22_X2 U2455 ( .A1(n419), .A2(n3180), .B1(n3179), .B2(n369), .ZN(n2622) );
  XOR2_X2 U2557 ( .A(a[16]), .B(n345), .Z(n3235) );
  NAND2_X4 U2577 ( .A1(n3242), .A2(n372), .ZN(n422) );
  NAND2_X4 U2580 ( .A1(n3243), .A2(n369), .ZN(n419) );
  NAND2_X1 U2585 ( .A1(n3801), .A2(n354), .ZN(n3696) );
  INV_X4 U2586 ( .A(a[24]), .ZN(n3801) );
  INV_X4 U2587 ( .A(a[2]), .ZN(n3572) );
  INV_X2 U2588 ( .A(n330), .ZN(n3289) );
  INV_X1 U2589 ( .A(n339), .ZN(n3286) );
  INV_X1 U2590 ( .A(n339), .ZN(n3717) );
  XNOR2_X1 U2591 ( .A(n465), .B(n327), .ZN(n3128) );
  AND2_X1 U2592 ( .A1(n465), .A2(n366), .ZN(n2093) );
  XNOR2_X1 U2593 ( .A(n465), .B(n333), .ZN(n3062) );
  XNOR2_X1 U2594 ( .A(n465), .B(n3425), .ZN(n3161) );
  XNOR2_X1 U2595 ( .A(n465), .B(n3681), .ZN(n3029) );
  XNOR2_X1 U2596 ( .A(n465), .B(n3571), .ZN(n2930) );
  XNOR2_X1 U2597 ( .A(n465), .B(n3640), .ZN(n3194) );
  XNOR2_X1 U2598 ( .A(n465), .B(n339), .ZN(n2996) );
  XNOR2_X1 U2599 ( .A(n465), .B(n354), .ZN(n2831) );
  XNOR2_X1 U2600 ( .A(n465), .B(n363), .ZN(n2732) );
  XNOR2_X1 U2601 ( .A(n465), .B(n3603), .ZN(n2963) );
  XNOR2_X1 U2602 ( .A(n465), .B(n360), .ZN(n2765) );
  XNOR2_X1 U2603 ( .A(n465), .B(n348), .ZN(n2897) );
  XNOR2_X1 U2604 ( .A(n465), .B(n351), .ZN(n2864) );
  XNOR2_X1 U2605 ( .A(n465), .B(n330), .ZN(n3095) );
  XNOR2_X1 U2606 ( .A(n465), .B(n366), .ZN(n2699) );
  XNOR2_X1 U2607 ( .A(n465), .B(n357), .ZN(n2798) );
  INV_X1 U2608 ( .A(n465), .ZN(n3812) );
  NAND2_X1 U2609 ( .A1(n3572), .A2(n321), .ZN(n3638) );
  XOR2_X1 U2610 ( .A(a[20]), .B(n351), .Z(n3233) );
  INV_X4 U2611 ( .A(a[14]), .ZN(n3410) );
  INV_X1 U2612 ( .A(a[30]), .ZN(n3724) );
  XOR2_X1 U2613 ( .A(a[6]), .B(n330), .Z(n3240) );
  INV_X1 U2614 ( .A(a[6]), .ZN(n3743) );
  INV_X1 U2615 ( .A(a[28]), .ZN(n3699) );
  NAND2_X1 U2616 ( .A1(a[16]), .A2(n342), .ZN(n3601) );
  INV_X1 U2617 ( .A(a[16]), .ZN(n3599) );
  INV_X2 U2618 ( .A(a[12]), .ZN(n3686) );
  AND2_X1 U2619 ( .A1(n465), .A2(a[0]), .ZN(product[0]) );
  OAI21_X1 U2620 ( .B1(a[0]), .B2(n3813), .A(n3640), .ZN(n2604) );
  INV_X1 U2621 ( .A(n511), .ZN(n2646) );
  XNOR2_X1 U2622 ( .A(n511), .B(n363), .ZN(n2710) );
  XNOR2_X1 U2623 ( .A(n511), .B(n360), .ZN(n2743) );
  XNOR2_X1 U2624 ( .A(n511), .B(n366), .ZN(n2677) );
  XNOR2_X1 U2625 ( .A(n511), .B(n3448), .ZN(n3007) );
  XNOR2_X1 U2626 ( .A(n511), .B(n351), .ZN(n2842) );
  XNOR2_X1 U2627 ( .A(n511), .B(n354), .ZN(n2809) );
  XNOR2_X1 U2628 ( .A(n511), .B(n357), .ZN(n2776) );
  XNOR2_X1 U2629 ( .A(n511), .B(n348), .ZN(n2875) );
  XNOR2_X1 U2630 ( .A(n511), .B(n339), .ZN(n2974) );
  XNOR2_X1 U2631 ( .A(n511), .B(n330), .ZN(n3073) );
  XNOR2_X1 U2632 ( .A(n511), .B(n342), .ZN(n2941) );
  XNOR2_X1 U2633 ( .A(n511), .B(n324), .ZN(n3139) );
  XNOR2_X1 U2634 ( .A(n511), .B(n327), .ZN(n3106) );
  XNOR2_X1 U2635 ( .A(n511), .B(n333), .ZN(n3040) );
  XNOR2_X1 U2636 ( .A(n511), .B(n3547), .ZN(n2908) );
  INV_X1 U2637 ( .A(n517), .ZN(n2643) );
  XNOR2_X1 U2638 ( .A(n517), .B(n366), .ZN(n2674) );
  XNOR2_X1 U2639 ( .A(n517), .B(n363), .ZN(n2707) );
  XNOR2_X1 U2640 ( .A(n517), .B(n357), .ZN(n2773) );
  XNOR2_X1 U2641 ( .A(n517), .B(n360), .ZN(n2740) );
  XNOR2_X1 U2642 ( .A(n517), .B(n339), .ZN(n2971) );
  XNOR2_X1 U2643 ( .A(n517), .B(n3571), .ZN(n2905) );
  XNOR2_X1 U2644 ( .A(n517), .B(n351), .ZN(n2839) );
  XNOR2_X1 U2645 ( .A(n517), .B(n354), .ZN(n2806) );
  XNOR2_X1 U2646 ( .A(n517), .B(n348), .ZN(n2872) );
  XNOR2_X1 U2647 ( .A(n517), .B(n327), .ZN(n3103) );
  XNOR2_X1 U2648 ( .A(n517), .B(n324), .ZN(n3136) );
  XNOR2_X1 U2649 ( .A(n517), .B(n3448), .ZN(n3004) );
  XNOR2_X1 U2650 ( .A(n517), .B(n330), .ZN(n3070) );
  XNOR2_X1 U2651 ( .A(n517), .B(n342), .ZN(n2938) );
  XNOR2_X1 U2652 ( .A(n517), .B(n333), .ZN(n3037) );
  INV_X1 U2653 ( .A(n515), .ZN(n2644) );
  XNOR2_X1 U2654 ( .A(n515), .B(n363), .ZN(n2708) );
  XNOR2_X1 U2655 ( .A(n515), .B(n366), .ZN(n2675) );
  XNOR2_X1 U2656 ( .A(n515), .B(n360), .ZN(n2741) );
  XNOR2_X1 U2657 ( .A(n515), .B(n357), .ZN(n2774) );
  XNOR2_X1 U2658 ( .A(n515), .B(n3571), .ZN(n2906) );
  XNOR2_X1 U2659 ( .A(n515), .B(n351), .ZN(n2840) );
  XNOR2_X1 U2660 ( .A(n515), .B(n339), .ZN(n2972) );
  XNOR2_X1 U2661 ( .A(n515), .B(n354), .ZN(n2807) );
  XNOR2_X1 U2662 ( .A(n515), .B(n330), .ZN(n3071) );
  XNOR2_X1 U2663 ( .A(n515), .B(n348), .ZN(n2873) );
  XNOR2_X1 U2664 ( .A(n515), .B(n327), .ZN(n3104) );
  XNOR2_X1 U2665 ( .A(n515), .B(n324), .ZN(n3137) );
  XNOR2_X1 U2666 ( .A(n515), .B(n342), .ZN(n2939) );
  XNOR2_X1 U2667 ( .A(n515), .B(n333), .ZN(n3038) );
  XNOR2_X1 U2668 ( .A(n515), .B(n3448), .ZN(n3005) );
  INV_X1 U2669 ( .A(n529), .ZN(n2637) );
  XNOR2_X1 U2670 ( .A(n529), .B(n366), .ZN(n2668) );
  XNOR2_X1 U2671 ( .A(n529), .B(n363), .ZN(n2701) );
  XNOR2_X1 U2672 ( .A(n529), .B(n360), .ZN(n2734) );
  XNOR2_X1 U2673 ( .A(n529), .B(n357), .ZN(n2767) );
  XNOR2_X1 U2674 ( .A(n529), .B(n348), .ZN(n2866) );
  XNOR2_X1 U2675 ( .A(n529), .B(n351), .ZN(n2833) );
  XNOR2_X1 U2676 ( .A(n529), .B(n354), .ZN(n2800) );
  XNOR2_X1 U2677 ( .A(n529), .B(n3571), .ZN(n2899) );
  XNOR2_X1 U2678 ( .A(n529), .B(n342), .ZN(n2932) );
  XNOR2_X1 U2679 ( .A(n529), .B(n3448), .ZN(n2998) );
  XNOR2_X1 U2680 ( .A(n529), .B(n339), .ZN(n2965) );
  XNOR2_X1 U2681 ( .A(n529), .B(n333), .ZN(n3031) );
  XNOR2_X1 U2682 ( .A(n529), .B(n327), .ZN(n3097) );
  XNOR2_X1 U2683 ( .A(n529), .B(n330), .ZN(n3064) );
  XNOR2_X1 U2684 ( .A(n529), .B(n324), .ZN(n3130) );
  INV_X1 U2685 ( .A(n523), .ZN(n2640) );
  XNOR2_X1 U2686 ( .A(n523), .B(n366), .ZN(n2671) );
  XNOR2_X1 U2687 ( .A(n523), .B(n363), .ZN(n2704) );
  XNOR2_X1 U2688 ( .A(n523), .B(n360), .ZN(n2737) );
  XNOR2_X1 U2689 ( .A(n523), .B(n354), .ZN(n2803) );
  XNOR2_X1 U2690 ( .A(n523), .B(n357), .ZN(n2770) );
  XNOR2_X1 U2691 ( .A(n523), .B(n351), .ZN(n2836) );
  XNOR2_X1 U2692 ( .A(n523), .B(n3547), .ZN(n2902) );
  XNOR2_X1 U2693 ( .A(n523), .B(n348), .ZN(n2869) );
  XNOR2_X1 U2694 ( .A(n523), .B(n339), .ZN(n2968) );
  XNOR2_X1 U2695 ( .A(n523), .B(n3550), .ZN(n3001) );
  XNOR2_X1 U2696 ( .A(n523), .B(n342), .ZN(n2935) );
  XNOR2_X1 U2697 ( .A(n523), .B(n324), .ZN(n3133) );
  XNOR2_X1 U2698 ( .A(n523), .B(n333), .ZN(n3034) );
  XNOR2_X1 U2699 ( .A(n523), .B(n330), .ZN(n3067) );
  XNOR2_X1 U2700 ( .A(n523), .B(n327), .ZN(n3100) );
  INV_X1 U2701 ( .A(n521), .ZN(n2641) );
  XNOR2_X1 U2702 ( .A(n521), .B(n366), .ZN(n2672) );
  XNOR2_X1 U2703 ( .A(n521), .B(n363), .ZN(n2705) );
  XNOR2_X1 U2704 ( .A(n521), .B(n357), .ZN(n2771) );
  XNOR2_X1 U2705 ( .A(n521), .B(n354), .ZN(n2804) );
  XNOR2_X1 U2706 ( .A(n521), .B(n351), .ZN(n2837) );
  XNOR2_X1 U2707 ( .A(n521), .B(n360), .ZN(n2738) );
  XNOR2_X1 U2708 ( .A(n521), .B(n3550), .ZN(n3002) );
  XNOR2_X1 U2709 ( .A(n521), .B(n348), .ZN(n2870) );
  XNOR2_X1 U2710 ( .A(n521), .B(n3571), .ZN(n2903) );
  XNOR2_X1 U2711 ( .A(n521), .B(n3603), .ZN(n2936) );
  XNOR2_X1 U2712 ( .A(n521), .B(n327), .ZN(n3101) );
  XNOR2_X1 U2713 ( .A(n521), .B(n330), .ZN(n3068) );
  XNOR2_X1 U2714 ( .A(n521), .B(n333), .ZN(n3035) );
  XNOR2_X1 U2715 ( .A(n521), .B(n324), .ZN(n3134) );
  XNOR2_X1 U2716 ( .A(n521), .B(n339), .ZN(n2969) );
  INV_X1 U2717 ( .A(n527), .ZN(n2638) );
  XNOR2_X1 U2718 ( .A(n527), .B(n366), .ZN(n2669) );
  XNOR2_X1 U2719 ( .A(n527), .B(n363), .ZN(n2702) );
  XNOR2_X1 U2720 ( .A(n527), .B(n360), .ZN(n2735) );
  XNOR2_X1 U2721 ( .A(n527), .B(n3775), .ZN(n2834) );
  XNOR2_X1 U2722 ( .A(n527), .B(n354), .ZN(n2801) );
  XNOR2_X1 U2723 ( .A(n527), .B(n357), .ZN(n2768) );
  XNOR2_X1 U2724 ( .A(n527), .B(n342), .ZN(n2933) );
  XNOR2_X1 U2725 ( .A(n527), .B(n3547), .ZN(n2900) );
  XNOR2_X1 U2726 ( .A(n527), .B(n3681), .ZN(n2999) );
  XNOR2_X1 U2727 ( .A(n527), .B(n348), .ZN(n2867) );
  XNOR2_X1 U2728 ( .A(n527), .B(n339), .ZN(n2966) );
  XNOR2_X1 U2729 ( .A(n527), .B(n327), .ZN(n3098) );
  XNOR2_X1 U2730 ( .A(n527), .B(n330), .ZN(n3065) );
  XNOR2_X1 U2731 ( .A(n527), .B(n324), .ZN(n3131) );
  XNOR2_X1 U2732 ( .A(n527), .B(n333), .ZN(n3032) );
  INV_X1 U2733 ( .A(n519), .ZN(n2642) );
  XNOR2_X1 U2734 ( .A(n519), .B(n366), .ZN(n2673) );
  XNOR2_X1 U2735 ( .A(n519), .B(n363), .ZN(n2706) );
  XNOR2_X1 U2736 ( .A(n519), .B(n357), .ZN(n2772) );
  XNOR2_X1 U2737 ( .A(n519), .B(n354), .ZN(n2805) );
  XNOR2_X1 U2738 ( .A(n519), .B(n351), .ZN(n2838) );
  XNOR2_X1 U2739 ( .A(n519), .B(n360), .ZN(n2739) );
  XNOR2_X1 U2740 ( .A(n519), .B(n3448), .ZN(n3003) );
  XNOR2_X1 U2741 ( .A(n519), .B(n348), .ZN(n2871) );
  XNOR2_X1 U2742 ( .A(n519), .B(n3571), .ZN(n2904) );
  XNOR2_X1 U2743 ( .A(n519), .B(n3603), .ZN(n2937) );
  XNOR2_X1 U2744 ( .A(n519), .B(n333), .ZN(n3036) );
  XNOR2_X1 U2745 ( .A(n519), .B(n324), .ZN(n3135) );
  XNOR2_X1 U2746 ( .A(n519), .B(n327), .ZN(n3102) );
  XNOR2_X1 U2747 ( .A(n519), .B(n339), .ZN(n2970) );
  XNOR2_X1 U2748 ( .A(n519), .B(n330), .ZN(n3069) );
  INV_X1 U2749 ( .A(n525), .ZN(n2639) );
  XNOR2_X1 U2750 ( .A(n525), .B(n366), .ZN(n2670) );
  XNOR2_X1 U2751 ( .A(n525), .B(n363), .ZN(n2703) );
  XNOR2_X1 U2752 ( .A(n525), .B(n360), .ZN(n2736) );
  XNOR2_X1 U2753 ( .A(n525), .B(n3775), .ZN(n2835) );
  XNOR2_X1 U2754 ( .A(n525), .B(n354), .ZN(n2802) );
  XNOR2_X1 U2755 ( .A(n525), .B(n3547), .ZN(n2901) );
  XNOR2_X1 U2756 ( .A(n525), .B(n357), .ZN(n2769) );
  XNOR2_X1 U2757 ( .A(n525), .B(n3550), .ZN(n3000) );
  XNOR2_X1 U2758 ( .A(n525), .B(n339), .ZN(n2967) );
  XNOR2_X1 U2759 ( .A(n525), .B(n342), .ZN(n2934) );
  XNOR2_X1 U2760 ( .A(n525), .B(n348), .ZN(n2868) );
  XNOR2_X1 U2761 ( .A(n525), .B(n324), .ZN(n3132) );
  XNOR2_X1 U2762 ( .A(n525), .B(n330), .ZN(n3066) );
  XNOR2_X1 U2763 ( .A(n525), .B(n333), .ZN(n3033) );
  XNOR2_X1 U2764 ( .A(n525), .B(n327), .ZN(n3099) );
  XNOR2_X1 U2765 ( .A(n469), .B(n333), .ZN(n3061) );
  XNOR2_X1 U2766 ( .A(n469), .B(n3425), .ZN(n3160) );
  XNOR2_X1 U2767 ( .A(n469), .B(n327), .ZN(n3127) );
  XNOR2_X1 U2768 ( .A(n469), .B(n3640), .ZN(n3193) );
  XNOR2_X1 U2769 ( .A(n469), .B(n3681), .ZN(n3028) );
  XNOR2_X1 U2770 ( .A(n469), .B(n339), .ZN(n2995) );
  INV_X1 U2771 ( .A(n469), .ZN(n2667) );
  XNOR2_X1 U2772 ( .A(n469), .B(n360), .ZN(n2764) );
  XNOR2_X1 U2773 ( .A(n469), .B(n342), .ZN(n2962) );
  XNOR2_X1 U2774 ( .A(n469), .B(n351), .ZN(n2863) );
  XNOR2_X1 U2775 ( .A(n469), .B(n354), .ZN(n2830) );
  XNOR2_X1 U2776 ( .A(n469), .B(n3547), .ZN(n2929) );
  XNOR2_X1 U2777 ( .A(n469), .B(n366), .ZN(n2698) );
  XNOR2_X1 U2778 ( .A(n469), .B(n348), .ZN(n2896) );
  XNOR2_X1 U2779 ( .A(n469), .B(n330), .ZN(n3094) );
  XNOR2_X1 U2780 ( .A(n469), .B(n357), .ZN(n2797) );
  XNOR2_X1 U2781 ( .A(n471), .B(n3425), .ZN(n3159) );
  XNOR2_X1 U2782 ( .A(n471), .B(n3640), .ZN(n3192) );
  XNOR2_X1 U2783 ( .A(n471), .B(n333), .ZN(n3060) );
  INV_X1 U2784 ( .A(n471), .ZN(n2666) );
  XNOR2_X1 U2785 ( .A(n471), .B(n327), .ZN(n3126) );
  XNOR2_X1 U2786 ( .A(n471), .B(n330), .ZN(n3093) );
  XNOR2_X1 U2787 ( .A(n471), .B(n3550), .ZN(n3027) );
  XNOR2_X1 U2788 ( .A(n471), .B(n339), .ZN(n2994) );
  XNOR2_X1 U2789 ( .A(n471), .B(n342), .ZN(n2961) );
  XNOR2_X1 U2790 ( .A(n471), .B(n351), .ZN(n2862) );
  XNOR2_X1 U2791 ( .A(n471), .B(n3547), .ZN(n2928) );
  XNOR2_X1 U2792 ( .A(n471), .B(n366), .ZN(n2697) );
  XNOR2_X1 U2793 ( .A(n471), .B(n348), .ZN(n2895) );
  XNOR2_X1 U2794 ( .A(n471), .B(n360), .ZN(n2763) );
  XNOR2_X1 U2795 ( .A(n471), .B(n357), .ZN(n2796) );
  XNOR2_X1 U2796 ( .A(n475), .B(n3640), .ZN(n3190) );
  INV_X1 U2797 ( .A(n475), .ZN(n2664) );
  XNOR2_X1 U2798 ( .A(n475), .B(n3425), .ZN(n3157) );
  XNOR2_X1 U2799 ( .A(n475), .B(n327), .ZN(n3124) );
  XNOR2_X1 U2800 ( .A(n475), .B(n330), .ZN(n3091) );
  XNOR2_X1 U2801 ( .A(n475), .B(n333), .ZN(n3058) );
  XNOR2_X1 U2802 ( .A(n475), .B(n354), .ZN(n2827) );
  XNOR2_X1 U2803 ( .A(n475), .B(n339), .ZN(n2992) );
  XNOR2_X1 U2804 ( .A(n475), .B(n357), .ZN(n2794) );
  XNOR2_X1 U2805 ( .A(n475), .B(n351), .ZN(n2860) );
  XNOR2_X1 U2806 ( .A(n475), .B(n360), .ZN(n2761) );
  XNOR2_X1 U2807 ( .A(n475), .B(n366), .ZN(n2695) );
  XNOR2_X1 U2808 ( .A(n475), .B(n348), .ZN(n2893) );
  XNOR2_X1 U2809 ( .A(n475), .B(n342), .ZN(n2959) );
  XNOR2_X1 U2810 ( .A(n475), .B(n3547), .ZN(n2926) );
  XNOR2_X1 U2811 ( .A(n475), .B(n363), .ZN(n2728) );
  XNOR2_X1 U2812 ( .A(n475), .B(n3448), .ZN(n3025) );
  INV_X1 U2813 ( .A(n513), .ZN(n2645) );
  XNOR2_X1 U2814 ( .A(n513), .B(n360), .ZN(n2742) );
  XNOR2_X1 U2815 ( .A(n513), .B(n363), .ZN(n2709) );
  XNOR2_X1 U2816 ( .A(n513), .B(n366), .ZN(n2676) );
  XNOR2_X1 U2817 ( .A(n513), .B(n354), .ZN(n2808) );
  XNOR2_X1 U2818 ( .A(n513), .B(n348), .ZN(n2874) );
  XNOR2_X1 U2819 ( .A(n513), .B(n357), .ZN(n2775) );
  XNOR2_X1 U2820 ( .A(n513), .B(n351), .ZN(n2841) );
  XNOR2_X1 U2821 ( .A(n513), .B(n333), .ZN(n3039) );
  XNOR2_X1 U2822 ( .A(n513), .B(n324), .ZN(n3138) );
  XNOR2_X1 U2823 ( .A(n513), .B(n342), .ZN(n2940) );
  XNOR2_X1 U2824 ( .A(n513), .B(n339), .ZN(n2973) );
  XNOR2_X1 U2825 ( .A(n513), .B(n330), .ZN(n3072) );
  XNOR2_X1 U2826 ( .A(n513), .B(n327), .ZN(n3105) );
  XNOR2_X1 U2827 ( .A(n513), .B(n345), .ZN(n2907) );
  XNOR2_X1 U2828 ( .A(n513), .B(n3448), .ZN(n3006) );
  XNOR2_X1 U2829 ( .A(n473), .B(n3425), .ZN(n3158) );
  XNOR2_X1 U2830 ( .A(n473), .B(n3640), .ZN(n3191) );
  INV_X1 U2831 ( .A(n473), .ZN(n2665) );
  XNOR2_X1 U2832 ( .A(n473), .B(n333), .ZN(n3059) );
  XNOR2_X1 U2833 ( .A(n473), .B(n327), .ZN(n3125) );
  XNOR2_X1 U2834 ( .A(n473), .B(n330), .ZN(n3092) );
  XNOR2_X1 U2835 ( .A(n473), .B(n351), .ZN(n2861) );
  XNOR2_X1 U2836 ( .A(n473), .B(n363), .ZN(n2729) );
  XNOR2_X1 U2837 ( .A(n473), .B(n3547), .ZN(n2927) );
  XNOR2_X1 U2838 ( .A(n473), .B(n339), .ZN(n2993) );
  XNOR2_X1 U2839 ( .A(n473), .B(n348), .ZN(n2894) );
  XNOR2_X1 U2840 ( .A(n473), .B(n342), .ZN(n2960) );
  XNOR2_X1 U2841 ( .A(n473), .B(n366), .ZN(n2696) );
  XNOR2_X1 U2842 ( .A(n473), .B(n360), .ZN(n2762) );
  XNOR2_X1 U2843 ( .A(n473), .B(n3448), .ZN(n3026) );
  XNOR2_X1 U2844 ( .A(n473), .B(n357), .ZN(n2795) );
  INV_X1 U2845 ( .A(n477), .ZN(n2663) );
  XNOR2_X1 U2846 ( .A(n477), .B(n330), .ZN(n3090) );
  XNOR2_X1 U2847 ( .A(n477), .B(n3640), .ZN(n3189) );
  XNOR2_X1 U2848 ( .A(n477), .B(n327), .ZN(n3123) );
  XNOR2_X1 U2849 ( .A(n477), .B(n324), .ZN(n3156) );
  XNOR2_X1 U2850 ( .A(n477), .B(n354), .ZN(n2826) );
  XNOR2_X1 U2851 ( .A(n477), .B(n357), .ZN(n2793) );
  XNOR2_X1 U2852 ( .A(n477), .B(n339), .ZN(n2991) );
  XNOR2_X1 U2853 ( .A(n477), .B(n342), .ZN(n2958) );
  XNOR2_X1 U2854 ( .A(n477), .B(n3448), .ZN(n3024) );
  XNOR2_X1 U2855 ( .A(n477), .B(n351), .ZN(n2859) );
  XNOR2_X1 U2856 ( .A(n477), .B(n360), .ZN(n2760) );
  XNOR2_X1 U2857 ( .A(n477), .B(n366), .ZN(n2694) );
  XNOR2_X1 U2858 ( .A(n477), .B(n3547), .ZN(n2925) );
  XNOR2_X1 U2859 ( .A(n477), .B(n348), .ZN(n2892) );
  XNOR2_X1 U2860 ( .A(n477), .B(n333), .ZN(n3057) );
  XNOR2_X1 U2861 ( .A(n477), .B(n363), .ZN(n2727) );
  INV_X1 U2862 ( .A(n483), .ZN(n2660) );
  XNOR2_X1 U2863 ( .A(n483), .B(n354), .ZN(n2823) );
  XNOR2_X1 U2864 ( .A(n483), .B(n363), .ZN(n2724) );
  XNOR2_X1 U2865 ( .A(n483), .B(n357), .ZN(n2790) );
  XNOR2_X1 U2866 ( .A(n483), .B(n324), .ZN(n3153) );
  XNOR2_X1 U2867 ( .A(n483), .B(n333), .ZN(n3054) );
  XNOR2_X1 U2868 ( .A(n483), .B(n366), .ZN(n2691) );
  XNOR2_X1 U2869 ( .A(n483), .B(n351), .ZN(n2856) );
  XNOR2_X1 U2870 ( .A(n483), .B(n342), .ZN(n2955) );
  XNOR2_X1 U2871 ( .A(n483), .B(n360), .ZN(n2757) );
  XNOR2_X1 U2872 ( .A(n483), .B(n348), .ZN(n2889) );
  XNOR2_X1 U2873 ( .A(n483), .B(n330), .ZN(n3087) );
  XNOR2_X1 U2874 ( .A(n483), .B(n327), .ZN(n3120) );
  XNOR2_X1 U2875 ( .A(n483), .B(n3547), .ZN(n2922) );
  XNOR2_X1 U2876 ( .A(n483), .B(n339), .ZN(n2988) );
  XNOR2_X1 U2877 ( .A(n483), .B(n3448), .ZN(n3021) );
  XNOR2_X1 U2878 ( .A(n479), .B(n3425), .ZN(n3155) );
  INV_X1 U2879 ( .A(n479), .ZN(n2662) );
  XNOR2_X1 U2880 ( .A(n479), .B(n357), .ZN(n2792) );
  XNOR2_X1 U2881 ( .A(n479), .B(n3547), .ZN(n2924) );
  XNOR2_X1 U2882 ( .A(n479), .B(n351), .ZN(n2858) );
  XNOR2_X1 U2883 ( .A(n479), .B(n3448), .ZN(n3023) );
  XNOR2_X1 U2884 ( .A(n479), .B(n330), .ZN(n3089) );
  XNOR2_X1 U2885 ( .A(n479), .B(n327), .ZN(n3122) );
  XNOR2_X1 U2886 ( .A(n479), .B(n342), .ZN(n2957) );
  XNOR2_X1 U2887 ( .A(n479), .B(n363), .ZN(n2726) );
  XNOR2_X1 U2888 ( .A(n479), .B(n339), .ZN(n2990) );
  XNOR2_X1 U2889 ( .A(n479), .B(n360), .ZN(n2759) );
  XNOR2_X1 U2890 ( .A(n479), .B(n366), .ZN(n2693) );
  XNOR2_X1 U2891 ( .A(n479), .B(n348), .ZN(n2891) );
  XNOR2_X1 U2892 ( .A(n479), .B(n333), .ZN(n3056) );
  INV_X1 U2893 ( .A(n481), .ZN(n2661) );
  XNOR2_X1 U2894 ( .A(n481), .B(n324), .ZN(n3154) );
  XNOR2_X1 U2895 ( .A(n481), .B(n333), .ZN(n3055) );
  XNOR2_X1 U2896 ( .A(n481), .B(n351), .ZN(n2857) );
  XNOR2_X1 U2897 ( .A(n481), .B(n357), .ZN(n2791) );
  XNOR2_X1 U2898 ( .A(n481), .B(n327), .ZN(n3121) );
  XNOR2_X1 U2899 ( .A(n481), .B(n366), .ZN(n2692) );
  XNOR2_X1 U2900 ( .A(n481), .B(n348), .ZN(n2890) );
  XNOR2_X1 U2901 ( .A(n481), .B(n363), .ZN(n2725) );
  XNOR2_X1 U2902 ( .A(n481), .B(n3448), .ZN(n3022) );
  XNOR2_X1 U2903 ( .A(n481), .B(n3547), .ZN(n2923) );
  XNOR2_X1 U2904 ( .A(n481), .B(n330), .ZN(n3088) );
  XNOR2_X1 U2905 ( .A(n481), .B(n342), .ZN(n2956) );
  XNOR2_X1 U2906 ( .A(n481), .B(n339), .ZN(n2989) );
  XNOR2_X1 U2907 ( .A(n481), .B(n360), .ZN(n2758) );
  INV_X1 U2908 ( .A(n485), .ZN(n2659) );
  XNOR2_X1 U2909 ( .A(n485), .B(n354), .ZN(n2822) );
  XNOR2_X1 U2910 ( .A(n485), .B(n363), .ZN(n2723) );
  XNOR2_X1 U2911 ( .A(n485), .B(n324), .ZN(n3152) );
  XNOR2_X1 U2912 ( .A(n485), .B(n357), .ZN(n2789) );
  XNOR2_X1 U2913 ( .A(n485), .B(n339), .ZN(n2987) );
  XNOR2_X1 U2914 ( .A(n485), .B(n330), .ZN(n3086) );
  XNOR2_X1 U2915 ( .A(n485), .B(n366), .ZN(n2690) );
  XNOR2_X1 U2916 ( .A(n485), .B(n333), .ZN(n3053) );
  XNOR2_X1 U2917 ( .A(n485), .B(n348), .ZN(n2888) );
  XNOR2_X1 U2918 ( .A(n485), .B(n351), .ZN(n2855) );
  XNOR2_X1 U2919 ( .A(n485), .B(n327), .ZN(n3119) );
  XNOR2_X1 U2920 ( .A(n485), .B(n360), .ZN(n2756) );
  XNOR2_X1 U2921 ( .A(n485), .B(n3547), .ZN(n2921) );
  XNOR2_X1 U2922 ( .A(n485), .B(n3448), .ZN(n3020) );
  XNOR2_X1 U2923 ( .A(n485), .B(n342), .ZN(n2954) );
  INV_X1 U2924 ( .A(n491), .ZN(n2656) );
  XNOR2_X1 U2925 ( .A(n491), .B(n333), .ZN(n3050) );
  XNOR2_X1 U2926 ( .A(n491), .B(n363), .ZN(n2720) );
  XNOR2_X1 U2927 ( .A(n491), .B(n366), .ZN(n2687) );
  XNOR2_X1 U2928 ( .A(n491), .B(n348), .ZN(n2885) );
  XNOR2_X1 U2929 ( .A(n491), .B(n357), .ZN(n2786) );
  XNOR2_X1 U2930 ( .A(n491), .B(n354), .ZN(n2819) );
  XNOR2_X1 U2931 ( .A(n491), .B(n327), .ZN(n3116) );
  XNOR2_X1 U2932 ( .A(n491), .B(n3448), .ZN(n3017) );
  XNOR2_X1 U2933 ( .A(n491), .B(n342), .ZN(n2951) );
  XNOR2_X1 U2934 ( .A(n491), .B(n3547), .ZN(n2918) );
  XNOR2_X1 U2935 ( .A(n491), .B(n330), .ZN(n3083) );
  XNOR2_X1 U2936 ( .A(n491), .B(n360), .ZN(n2753) );
  XNOR2_X1 U2937 ( .A(n491), .B(n339), .ZN(n2984) );
  XNOR2_X1 U2938 ( .A(n491), .B(n351), .ZN(n2852) );
  XNOR2_X1 U2939 ( .A(n491), .B(n324), .ZN(n3149) );
  INV_X1 U2940 ( .A(n487), .ZN(n2658) );
  XNOR2_X1 U2941 ( .A(n487), .B(n366), .ZN(n2689) );
  XNOR2_X1 U2942 ( .A(n487), .B(n324), .ZN(n3151) );
  XNOR2_X1 U2943 ( .A(n487), .B(n330), .ZN(n3085) );
  XNOR2_X1 U2944 ( .A(n487), .B(n339), .ZN(n2986) );
  XNOR2_X1 U2945 ( .A(n487), .B(n357), .ZN(n2788) );
  XNOR2_X1 U2946 ( .A(n487), .B(n327), .ZN(n3118) );
  XNOR2_X1 U2947 ( .A(n487), .B(n351), .ZN(n2854) );
  XNOR2_X1 U2948 ( .A(n487), .B(n360), .ZN(n2755) );
  XNOR2_X1 U2949 ( .A(n487), .B(n363), .ZN(n2722) );
  XNOR2_X1 U2950 ( .A(n487), .B(n345), .ZN(n2920) );
  XNOR2_X1 U2951 ( .A(n487), .B(n348), .ZN(n2887) );
  XNOR2_X1 U2952 ( .A(n487), .B(n333), .ZN(n3052) );
  XNOR2_X1 U2953 ( .A(n487), .B(n3448), .ZN(n3019) );
  XNOR2_X1 U2954 ( .A(n487), .B(n342), .ZN(n2953) );
  INV_X1 U2955 ( .A(n489), .ZN(n2657) );
  XNOR2_X1 U2956 ( .A(n489), .B(n330), .ZN(n3084) );
  XNOR2_X1 U2957 ( .A(n489), .B(n357), .ZN(n2787) );
  XNOR2_X1 U2958 ( .A(n489), .B(n333), .ZN(n3051) );
  XNOR2_X1 U2959 ( .A(n489), .B(n366), .ZN(n2688) );
  XNOR2_X1 U2960 ( .A(n489), .B(n363), .ZN(n2721) );
  XNOR2_X1 U2961 ( .A(n489), .B(n342), .ZN(n2952) );
  XNOR2_X1 U2962 ( .A(n489), .B(n327), .ZN(n3117) );
  XNOR2_X1 U2963 ( .A(n489), .B(n348), .ZN(n2886) );
  XNOR2_X1 U2964 ( .A(n489), .B(n360), .ZN(n2754) );
  XNOR2_X1 U2965 ( .A(n489), .B(n3448), .ZN(n3018) );
  XNOR2_X1 U2966 ( .A(n489), .B(n3547), .ZN(n2919) );
  XNOR2_X1 U2967 ( .A(n489), .B(n339), .ZN(n2985) );
  XNOR2_X1 U2968 ( .A(n489), .B(n351), .ZN(n2853) );
  XNOR2_X1 U2969 ( .A(n489), .B(n324), .ZN(n3150) );
  INV_X1 U2970 ( .A(n493), .ZN(n2655) );
  XNOR2_X1 U2971 ( .A(n493), .B(n366), .ZN(n2686) );
  XNOR2_X1 U2972 ( .A(n493), .B(n363), .ZN(n2719) );
  XNOR2_X1 U2973 ( .A(n493), .B(n345), .ZN(n2917) );
  XNOR2_X1 U2974 ( .A(n493), .B(n333), .ZN(n3049) );
  XNOR2_X1 U2975 ( .A(n493), .B(n324), .ZN(n3148) );
  XNOR2_X1 U2976 ( .A(n493), .B(n3550), .ZN(n3016) );
  XNOR2_X1 U2977 ( .A(n493), .B(n348), .ZN(n2884) );
  XNOR2_X1 U2978 ( .A(n493), .B(n354), .ZN(n2818) );
  XNOR2_X1 U2979 ( .A(n493), .B(n342), .ZN(n2950) );
  XNOR2_X1 U2980 ( .A(n493), .B(n357), .ZN(n2785) );
  XNOR2_X1 U2981 ( .A(n493), .B(n327), .ZN(n3115) );
  XNOR2_X1 U2982 ( .A(n493), .B(n360), .ZN(n2752) );
  XNOR2_X1 U2983 ( .A(n493), .B(n339), .ZN(n2983) );
  XNOR2_X1 U2984 ( .A(n493), .B(n330), .ZN(n3082) );
  XNOR2_X1 U2985 ( .A(n493), .B(n351), .ZN(n2851) );
  INV_X1 U2986 ( .A(n499), .ZN(n2652) );
  XNOR2_X1 U2987 ( .A(n499), .B(n366), .ZN(n2683) );
  XNOR2_X1 U2988 ( .A(n499), .B(n363), .ZN(n2716) );
  XNOR2_X1 U2989 ( .A(n499), .B(n357), .ZN(n2782) );
  XNOR2_X1 U2990 ( .A(n499), .B(n360), .ZN(n2749) );
  XNOR2_X1 U2991 ( .A(n499), .B(n354), .ZN(n2815) );
  XNOR2_X1 U2992 ( .A(n499), .B(n3547), .ZN(n2914) );
  XNOR2_X1 U2993 ( .A(n499), .B(n3448), .ZN(n3013) );
  XNOR2_X1 U2994 ( .A(n499), .B(n342), .ZN(n2947) );
  XNOR2_X1 U2995 ( .A(n499), .B(n351), .ZN(n2848) );
  XNOR2_X1 U2996 ( .A(n499), .B(n330), .ZN(n3079) );
  XNOR2_X1 U2997 ( .A(n499), .B(n324), .ZN(n3145) );
  XNOR2_X1 U2998 ( .A(n499), .B(n327), .ZN(n3112) );
  XNOR2_X1 U2999 ( .A(n499), .B(n348), .ZN(n2881) );
  XNOR2_X1 U3000 ( .A(n499), .B(n333), .ZN(n3046) );
  INV_X1 U3001 ( .A(n495), .ZN(n2654) );
  XNOR2_X1 U3002 ( .A(n495), .B(n366), .ZN(n2685) );
  XNOR2_X1 U3003 ( .A(n495), .B(n363), .ZN(n2718) );
  XNOR2_X1 U3004 ( .A(n495), .B(n360), .ZN(n2751) );
  XNOR2_X1 U3005 ( .A(n495), .B(n354), .ZN(n2817) );
  XNOR2_X1 U3006 ( .A(n495), .B(n339), .ZN(n2982) );
  XNOR2_X1 U3007 ( .A(n495), .B(n3547), .ZN(n2916) );
  XNOR2_X1 U3008 ( .A(n495), .B(n333), .ZN(n3048) );
  XNOR2_X1 U3009 ( .A(n495), .B(n324), .ZN(n3147) );
  XNOR2_X1 U3010 ( .A(n495), .B(n351), .ZN(n2850) );
  XNOR2_X1 U3011 ( .A(n495), .B(n330), .ZN(n3081) );
  XNOR2_X1 U3012 ( .A(n495), .B(n3448), .ZN(n3015) );
  XNOR2_X1 U3013 ( .A(n495), .B(n348), .ZN(n2883) );
  XNOR2_X1 U3014 ( .A(n495), .B(n357), .ZN(n2784) );
  XNOR2_X1 U3015 ( .A(n495), .B(n327), .ZN(n3114) );
  XNOR2_X1 U3016 ( .A(n495), .B(n342), .ZN(n2949) );
  INV_X1 U3017 ( .A(n497), .ZN(n2653) );
  XNOR2_X1 U3018 ( .A(n497), .B(n366), .ZN(n2684) );
  XNOR2_X1 U3019 ( .A(n497), .B(n354), .ZN(n2816) );
  XNOR2_X1 U3020 ( .A(n497), .B(n363), .ZN(n2717) );
  XNOR2_X1 U3021 ( .A(n497), .B(n360), .ZN(n2750) );
  XNOR2_X1 U3022 ( .A(n497), .B(n324), .ZN(n3146) );
  XNOR2_X1 U3023 ( .A(n497), .B(n3547), .ZN(n2915) );
  XNOR2_X1 U3024 ( .A(n497), .B(n351), .ZN(n2849) );
  XNOR2_X1 U3025 ( .A(n497), .B(n357), .ZN(n2783) );
  XNOR2_X1 U3026 ( .A(n497), .B(n330), .ZN(n3080) );
  XNOR2_X1 U3027 ( .A(n497), .B(n3448), .ZN(n3014) );
  XNOR2_X1 U3028 ( .A(n497), .B(n348), .ZN(n2882) );
  XNOR2_X1 U3029 ( .A(n497), .B(n342), .ZN(n2948) );
  XNOR2_X1 U3030 ( .A(n497), .B(n333), .ZN(n3047) );
  XNOR2_X1 U3031 ( .A(n497), .B(n327), .ZN(n3113) );
  INV_X1 U3032 ( .A(n501), .ZN(n2651) );
  XNOR2_X1 U3033 ( .A(n501), .B(n366), .ZN(n2682) );
  XNOR2_X1 U3034 ( .A(n501), .B(n360), .ZN(n2748) );
  XNOR2_X1 U3035 ( .A(n501), .B(n357), .ZN(n2781) );
  XNOR2_X1 U3036 ( .A(n501), .B(n363), .ZN(n2715) );
  XNOR2_X1 U3037 ( .A(n501), .B(n351), .ZN(n2847) );
  XNOR2_X1 U3038 ( .A(n501), .B(n327), .ZN(n3111) );
  XNOR2_X1 U3039 ( .A(n501), .B(n339), .ZN(n2979) );
  XNOR2_X1 U3040 ( .A(n501), .B(n342), .ZN(n2946) );
  XNOR2_X1 U3041 ( .A(n501), .B(n330), .ZN(n3078) );
  XNOR2_X1 U3042 ( .A(n501), .B(n354), .ZN(n2814) );
  XNOR2_X1 U3043 ( .A(n501), .B(n3448), .ZN(n3012) );
  XNOR2_X1 U3044 ( .A(n501), .B(n3547), .ZN(n2913) );
  XNOR2_X1 U3045 ( .A(n501), .B(n324), .ZN(n3144) );
  XNOR2_X1 U3046 ( .A(n501), .B(n333), .ZN(n3045) );
  XNOR2_X1 U3047 ( .A(n501), .B(n348), .ZN(n2880) );
  INV_X1 U3048 ( .A(n505), .ZN(n2649) );
  XNOR2_X1 U3049 ( .A(n505), .B(n366), .ZN(n2680) );
  XNOR2_X1 U3050 ( .A(n505), .B(n3550), .ZN(n3010) );
  XNOR2_X1 U3051 ( .A(n505), .B(n363), .ZN(n2713) );
  XNOR2_X1 U3052 ( .A(n505), .B(n360), .ZN(n2746) );
  XNOR2_X1 U3053 ( .A(n505), .B(n354), .ZN(n2812) );
  XNOR2_X1 U3054 ( .A(n505), .B(n351), .ZN(n2845) );
  XNOR2_X1 U3055 ( .A(n505), .B(n357), .ZN(n2779) );
  XNOR2_X1 U3056 ( .A(n505), .B(n339), .ZN(n2977) );
  XNOR2_X1 U3057 ( .A(n505), .B(n330), .ZN(n3076) );
  XNOR2_X1 U3058 ( .A(n505), .B(n3547), .ZN(n2911) );
  XNOR2_X1 U3059 ( .A(n505), .B(n324), .ZN(n3142) );
  XNOR2_X1 U3060 ( .A(n505), .B(n327), .ZN(n3109) );
  XNOR2_X1 U3061 ( .A(n505), .B(n333), .ZN(n3043) );
  XNOR2_X1 U3062 ( .A(n505), .B(n342), .ZN(n2944) );
  INV_X1 U3063 ( .A(n503), .ZN(n2650) );
  XNOR2_X1 U3064 ( .A(n503), .B(n363), .ZN(n2714) );
  XNOR2_X1 U3065 ( .A(n503), .B(n366), .ZN(n2681) );
  XNOR2_X1 U3066 ( .A(n503), .B(n360), .ZN(n2747) );
  XNOR2_X1 U3067 ( .A(n503), .B(n354), .ZN(n2813) );
  XNOR2_X1 U3068 ( .A(n503), .B(n351), .ZN(n2846) );
  XNOR2_X1 U3069 ( .A(n503), .B(n357), .ZN(n2780) );
  XNOR2_X1 U3070 ( .A(n503), .B(n327), .ZN(n3110) );
  XNOR2_X1 U3071 ( .A(n503), .B(n333), .ZN(n3044) );
  XNOR2_X1 U3072 ( .A(n503), .B(n330), .ZN(n3077) );
  XNOR2_X1 U3073 ( .A(n503), .B(n339), .ZN(n2978) );
  XNOR2_X1 U3074 ( .A(n503), .B(n324), .ZN(n3143) );
  XNOR2_X1 U3075 ( .A(n503), .B(n3448), .ZN(n3011) );
  XNOR2_X1 U3076 ( .A(n503), .B(n342), .ZN(n2945) );
  XNOR2_X1 U3077 ( .A(n503), .B(n345), .ZN(n2912) );
  INV_X1 U3078 ( .A(n507), .ZN(n2648) );
  XNOR2_X1 U3079 ( .A(n507), .B(n366), .ZN(n2679) );
  XNOR2_X1 U3080 ( .A(n507), .B(n363), .ZN(n2712) );
  XNOR2_X1 U3081 ( .A(n507), .B(n360), .ZN(n2745) );
  XNOR2_X1 U3082 ( .A(n507), .B(n357), .ZN(n2778) );
  XNOR2_X1 U3083 ( .A(n507), .B(n354), .ZN(n2811) );
  XNOR2_X1 U3084 ( .A(n507), .B(n3550), .ZN(n3009) );
  XNOR2_X1 U3085 ( .A(n507), .B(n339), .ZN(n2976) );
  XNOR2_X1 U3086 ( .A(n507), .B(n351), .ZN(n2844) );
  XNOR2_X1 U3087 ( .A(n507), .B(n324), .ZN(n3141) );
  XNOR2_X1 U3088 ( .A(n507), .B(n330), .ZN(n3075) );
  XNOR2_X1 U3089 ( .A(n507), .B(n348), .ZN(n2877) );
  XNOR2_X1 U3090 ( .A(n507), .B(n333), .ZN(n3042) );
  XNOR2_X1 U3091 ( .A(n507), .B(n327), .ZN(n3108) );
  XNOR2_X1 U3092 ( .A(n507), .B(n3547), .ZN(n2910) );
  XNOR2_X1 U3093 ( .A(n507), .B(n342), .ZN(n2943) );
  INV_X1 U3094 ( .A(n509), .ZN(n2647) );
  XNOR2_X1 U3095 ( .A(n509), .B(n363), .ZN(n2711) );
  XNOR2_X1 U3096 ( .A(n509), .B(n366), .ZN(n2678) );
  XNOR2_X1 U3097 ( .A(n509), .B(n360), .ZN(n2744) );
  XNOR2_X1 U3098 ( .A(n509), .B(n330), .ZN(n3074) );
  XNOR2_X1 U3099 ( .A(n509), .B(n354), .ZN(n2810) );
  XNOR2_X1 U3100 ( .A(n509), .B(n357), .ZN(n2777) );
  XNOR2_X1 U3101 ( .A(n509), .B(n351), .ZN(n2843) );
  XNOR2_X1 U3102 ( .A(n509), .B(n3448), .ZN(n3008) );
  XNOR2_X1 U3103 ( .A(n509), .B(n339), .ZN(n2975) );
  XNOR2_X1 U3104 ( .A(n509), .B(n324), .ZN(n3140) );
  XNOR2_X1 U3105 ( .A(n509), .B(n333), .ZN(n3041) );
  XNOR2_X1 U3106 ( .A(n509), .B(n348), .ZN(n2876) );
  XNOR2_X1 U3107 ( .A(n509), .B(n345), .ZN(n2909) );
  XNOR2_X1 U3108 ( .A(n509), .B(n327), .ZN(n3107) );
  XNOR2_X1 U3109 ( .A(n509), .B(n342), .ZN(n2942) );
  NAND2_X2 U3110 ( .A1(n3606), .A2(n345), .ZN(n3609) );
  XOR2_X1 U3111 ( .A(n3583), .B(n3290), .Z(n3241) );
  INV_X4 U3112 ( .A(n327), .ZN(n3290) );
  NAND3_X1 U3113 ( .A1(n3713), .A2(n3715), .A3(n3714), .ZN(n3409) );
  NAND3_X1 U3114 ( .A1(n3713), .A2(n3715), .A3(n3714), .ZN(n1518) );
  OAI22_X2 U3115 ( .A1(n3723), .A2(n3130), .B1(n372), .B2(n3291), .ZN(n2571)
         );
  NOR2_X1 U3116 ( .A1(n727), .A2(n688), .ZN(n3411) );
  NOR2_X1 U3117 ( .A1(n727), .A2(n688), .ZN(n686) );
  NOR2_X2 U3118 ( .A1(n1519), .A2(n1550), .ZN(n3754) );
  INV_X1 U3119 ( .A(n3734), .ZN(n3735) );
  XNOR2_X1 U3120 ( .A(n1552), .B(n1523), .ZN(n3675) );
  NAND2_X1 U3121 ( .A1(n3410), .A2(n339), .ZN(n3718) );
  XNOR2_X1 U3122 ( .A(n3801), .B(n357), .ZN(n3231) );
  XNOR2_X1 U3123 ( .A(n3615), .B(n360), .ZN(n3230) );
  INV_X4 U3124 ( .A(a[26]), .ZN(n3615) );
  NAND2_X1 U3125 ( .A1(n752), .A2(n729), .ZN(n727) );
  XOR2_X1 U3126 ( .A(n2156), .B(n1580), .Z(n3412) );
  XOR2_X1 U3127 ( .A(n2412), .B(n3412), .Z(n1579) );
  NAND2_X1 U3128 ( .A1(n2412), .A2(n2156), .ZN(n3413) );
  NAND2_X1 U3129 ( .A1(n2412), .A2(n1580), .ZN(n3414) );
  NAND2_X1 U3130 ( .A1(n2156), .A2(n1580), .ZN(n3415) );
  NAND3_X1 U3131 ( .A1(n3413), .A2(n3415), .A3(n3414), .ZN(n1578) );
  XOR2_X1 U3132 ( .A(n1566), .B(n1568), .Z(n3416) );
  XOR2_X1 U3133 ( .A(n3416), .B(n1564), .Z(n1529) );
  XOR2_X1 U3134 ( .A(n1558), .B(n1527), .Z(n3417) );
  XOR2_X1 U3135 ( .A(n3417), .B(n1529), .Z(n1523) );
  NAND2_X1 U3136 ( .A1(n1566), .A2(n1568), .ZN(n3418) );
  NAND2_X1 U3137 ( .A1(n1566), .A2(n1564), .ZN(n3419) );
  NAND2_X1 U3138 ( .A1(n1568), .A2(n1564), .ZN(n3420) );
  NAND3_X1 U3139 ( .A1(n3418), .A2(n3419), .A3(n3420), .ZN(n1528) );
  NAND2_X1 U3140 ( .A1(n1558), .A2(n1527), .ZN(n3421) );
  NAND2_X1 U3141 ( .A1(n1558), .A2(n1529), .ZN(n3422) );
  NAND2_X1 U3142 ( .A1(n1527), .A2(n1529), .ZN(n3423) );
  NAND3_X1 U3143 ( .A1(n3421), .A2(n3422), .A3(n3423), .ZN(n1522) );
  INV_X1 U3144 ( .A(n1548), .ZN(n1580) );
  INV_X4 U3145 ( .A(n324), .ZN(n3424) );
  INV_X2 U3146 ( .A(n3424), .ZN(n3425) );
  NAND2_X2 U3147 ( .A1(n3242), .A2(n372), .ZN(n3723) );
  INV_X1 U3148 ( .A(n753), .ZN(n751) );
  OAI22_X1 U3149 ( .A1(n446), .A2(n2895), .B1(n2894), .B2(n3729), .ZN(n2328)
         );
  OAI22_X1 U3150 ( .A1(n446), .A2(n2897), .B1(n2896), .B2(n3729), .ZN(n2330)
         );
  OAI22_X1 U3151 ( .A1(n446), .A2(n2892), .B1(n2891), .B2(n3728), .ZN(n2325)
         );
  OAI22_X1 U3152 ( .A1(n446), .A2(n2884), .B1(n2883), .B2(n3728), .ZN(n2317)
         );
  OAI22_X1 U3153 ( .A1(n446), .A2(n2882), .B1(n2881), .B2(n3728), .ZN(n2315)
         );
  AND2_X2 U3154 ( .A1(n3234), .A2(n3727), .ZN(n3803) );
  XOR2_X1 U3155 ( .A(n2387), .B(n2515), .Z(n3426) );
  XOR2_X1 U3156 ( .A(n3426), .B(n2419), .Z(n1766) );
  XOR2_X1 U3157 ( .A(n1793), .B(n1768), .Z(n3427) );
  XOR2_X1 U3158 ( .A(n3427), .B(n1766), .Z(n1760) );
  NAND2_X1 U3159 ( .A1(n2387), .A2(n2515), .ZN(n3428) );
  NAND2_X1 U3160 ( .A1(n2387), .A2(n2419), .ZN(n3429) );
  NAND2_X1 U3161 ( .A1(n2515), .A2(n2419), .ZN(n3430) );
  NAND3_X1 U3162 ( .A1(n3428), .A2(n3429), .A3(n3430), .ZN(n1765) );
  NAND2_X1 U3163 ( .A1(n1793), .A2(n1768), .ZN(n3431) );
  NAND2_X1 U3164 ( .A1(n1793), .A2(n1766), .ZN(n3432) );
  NAND2_X1 U3165 ( .A1(n1768), .A2(n1766), .ZN(n3433) );
  NAND3_X1 U3166 ( .A1(n3431), .A2(n3432), .A3(n3433), .ZN(n1759) );
  XOR2_X1 U3167 ( .A(n1751), .B(n1728), .Z(n3434) );
  XOR2_X1 U3168 ( .A(n1726), .B(n3434), .Z(n1724) );
  NAND2_X1 U3169 ( .A1(n1726), .A2(n1751), .ZN(n3435) );
  NAND2_X1 U3170 ( .A1(n1726), .A2(n1728), .ZN(n3436) );
  NAND2_X1 U3171 ( .A1(n1751), .A2(n1728), .ZN(n3437) );
  NAND3_X1 U3172 ( .A1(n3435), .A2(n3437), .A3(n3436), .ZN(n1723) );
  XOR2_X1 U3173 ( .A(a[12]), .B(n339), .Z(n3237) );
  XOR2_X1 U3174 ( .A(a[8]), .B(n333), .Z(n3239) );
  NOR2_X1 U3175 ( .A1(n861), .A2(n864), .ZN(n3438) );
  NOR2_X1 U3176 ( .A1(n861), .A2(n864), .ZN(n859) );
  INV_X1 U3177 ( .A(n3494), .ZN(n3439) );
  AND2_X2 U3178 ( .A1(n3230), .A2(n408), .ZN(n3808) );
  NAND2_X2 U3179 ( .A1(n1519), .A2(n1550), .ZN(n794) );
  XOR2_X1 U3180 ( .A(a[28]), .B(n363), .Z(n3229) );
  INV_X1 U3181 ( .A(n3445), .ZN(n3790) );
  INV_X1 U3182 ( .A(n3445), .ZN(n3676) );
  BUF_X1 U3183 ( .A(n1520), .Z(n3440) );
  NAND2_X2 U3184 ( .A1(n3617), .A2(n3618), .ZN(n3792) );
  NAND2_X2 U3185 ( .A1(n3228), .A2(n3641), .ZN(n3457) );
  NOR2_X1 U3186 ( .A1(n819), .A2(n824), .ZN(n817) );
  AND2_X2 U3187 ( .A1(n3231), .A2(n405), .ZN(n3580) );
  BUF_X1 U3188 ( .A(n3778), .Z(n3441) );
  OAI21_X1 U3189 ( .B1(n660), .B2(n664), .A(n661), .ZN(n659) );
  AOI21_X2 U3190 ( .B1(n612), .B2(n981), .A(n607), .ZN(n605) );
  AOI21_X1 U3191 ( .B1(n844), .B2(n852), .A(n845), .ZN(n3442) );
  AOI21_X1 U3192 ( .B1(n844), .B2(n852), .A(n845), .ZN(n843) );
  INV_X1 U3193 ( .A(n711), .ZN(n709) );
  NOR2_X1 U3194 ( .A1(n692), .A2(n711), .ZN(n690) );
  INV_X2 U3195 ( .A(n3812), .ZN(n3443) );
  INV_X8 U3196 ( .A(n3443), .ZN(n3444) );
  AND2_X2 U3197 ( .A1(n3745), .A2(n3746), .ZN(n3445) );
  OAI22_X1 U3198 ( .A1(n3705), .A2(n2784), .B1(n2783), .B2(n3581), .ZN(n2214)
         );
  INV_X8 U3199 ( .A(n3579), .ZN(n3705) );
  NAND2_X1 U3200 ( .A1(n3686), .A2(n336), .ZN(n3689) );
  BUF_X1 U3201 ( .A(n861), .Z(n3446) );
  XNOR2_X1 U3202 ( .A(n3447), .B(n1451), .ZN(n1443) );
  XNOR2_X1 U3203 ( .A(n1449), .B(n1457), .ZN(n3447) );
  BUF_X8 U3204 ( .A(n336), .Z(n3448) );
  OAI22_X1 U3205 ( .A1(n3723), .A2(n3291), .B1(n3162), .B2(n3573), .ZN(n2075)
         );
  OAI22_X1 U3206 ( .A1(n3723), .A2(n3160), .B1(n3159), .B2(n3573), .ZN(n2601)
         );
  OAI22_X1 U3207 ( .A1(n3723), .A2(n3157), .B1(n3156), .B2(n3573), .ZN(n2598)
         );
  OAI22_X1 U3208 ( .A1(n3723), .A2(n3152), .B1(n3151), .B2(n3573), .ZN(n2593)
         );
  OAI22_X1 U3209 ( .A1(n3723), .A2(n3148), .B1(n3147), .B2(n3573), .ZN(n2589)
         );
  OAI22_X1 U3210 ( .A1(n3723), .A2(n3133), .B1(n3132), .B2(n3573), .ZN(n2574)
         );
  OAI22_X1 U3211 ( .A1(n3723), .A2(n3151), .B1(n3150), .B2(n3573), .ZN(n2592)
         );
  OAI22_X1 U3212 ( .A1(n3723), .A2(n3138), .B1(n3137), .B2(n3573), .ZN(n2579)
         );
  OAI22_X1 U3213 ( .A1(n3723), .A2(n3140), .B1(n3139), .B2(n3573), .ZN(n2581)
         );
  NOR2_X1 U3214 ( .A1(n1820), .A2(n1841), .ZN(n3475) );
  OAI22_X1 U3215 ( .A1(n422), .A2(n3158), .B1(n3157), .B2(n3573), .ZN(n2599)
         );
  OAI22_X1 U3216 ( .A1(n422), .A2(n3147), .B1(n3146), .B2(n3573), .ZN(n2588)
         );
  OAI22_X1 U3217 ( .A1(n422), .A2(n3155), .B1(n3154), .B2(n3573), .ZN(n2596)
         );
  OAI22_X1 U3218 ( .A1(n422), .A2(n3154), .B1(n3153), .B2(n3573), .ZN(n2595)
         );
  OAI22_X1 U3219 ( .A1(n422), .A2(n3136), .B1(n3135), .B2(n3573), .ZN(n2577)
         );
  OAI22_X1 U3220 ( .A1(n422), .A2(n3135), .B1(n3134), .B2(n3573), .ZN(n2576)
         );
  OAI22_X1 U3221 ( .A1(n422), .A2(n3144), .B1(n3143), .B2(n3573), .ZN(n2585)
         );
  OAI22_X1 U3222 ( .A1(n422), .A2(n3139), .B1(n3138), .B2(n3573), .ZN(n2580)
         );
  OAI22_X1 U3223 ( .A1(n422), .A2(n3141), .B1(n3140), .B2(n3573), .ZN(n2582)
         );
  OAI22_X1 U3224 ( .A1(n422), .A2(n3150), .B1(n3149), .B2(n372), .ZN(n2591) );
  NAND2_X1 U3225 ( .A1(n994), .A2(n705), .ZN(n548) );
  NAND2_X2 U3226 ( .A1(n694), .A2(n994), .ZN(n692) );
  NAND2_X1 U3227 ( .A1(n1201), .A2(n1218), .ZN(n705) );
  NOR2_X1 U3228 ( .A1(n1201), .A2(n1218), .ZN(n704) );
  XOR2_X1 U3229 ( .A(n1590), .B(n1588), .Z(n3449) );
  XOR2_X1 U3230 ( .A(n3449), .B(n1615), .Z(n1584) );
  XOR2_X1 U3231 ( .A(n1613), .B(n1586), .Z(n3450) );
  XOR2_X1 U3232 ( .A(n3450), .B(n1584), .Z(n1582) );
  NAND2_X1 U3233 ( .A1(n1590), .A2(n1588), .ZN(n3451) );
  NAND2_X1 U3234 ( .A1(n1590), .A2(n1615), .ZN(n3452) );
  NAND2_X1 U3235 ( .A1(n1588), .A2(n1615), .ZN(n3453) );
  NAND3_X1 U3236 ( .A1(n3451), .A2(n3452), .A3(n3453), .ZN(n1583) );
  NAND2_X1 U3237 ( .A1(n1613), .A2(n1586), .ZN(n3454) );
  NAND2_X1 U3238 ( .A1(n1613), .A2(n1584), .ZN(n3455) );
  NAND2_X1 U3239 ( .A1(n1586), .A2(n1584), .ZN(n3456) );
  NAND3_X1 U3240 ( .A1(n3454), .A2(n3455), .A3(n3456), .ZN(n1581) );
  INV_X1 U3241 ( .A(n399), .ZN(n3611) );
  OAI22_X1 U3242 ( .A1(n3620), .A2(n3065), .B1(n3064), .B2(n3679), .ZN(n2504)
         );
  XNOR2_X2 U3243 ( .A(a[0]), .B(n3637), .ZN(n3243) );
  INV_X4 U3244 ( .A(n321), .ZN(n3637) );
  AND2_X1 U3245 ( .A1(n3238), .A2(n3588), .ZN(n3732) );
  INV_X2 U3246 ( .A(n3806), .ZN(n3788) );
  NAND2_X4 U3247 ( .A1(n3228), .A2(n3641), .ZN(n3458) );
  XOR2_X2 U3248 ( .A(a[30]), .B(n366), .Z(n3228) );
  INV_X2 U3249 ( .A(n3792), .ZN(n3741) );
  INV_X2 U3250 ( .A(n3792), .ZN(n3742) );
  AOI21_X2 U3251 ( .B1(n3604), .B2(n838), .A(n833), .ZN(n831) );
  XOR2_X1 U3252 ( .A(n1384), .B(n1361), .Z(n3459) );
  XOR2_X1 U3253 ( .A(n1359), .B(n3459), .Z(n1355) );
  NAND2_X1 U3254 ( .A1(n1359), .A2(n1384), .ZN(n3460) );
  NAND2_X1 U3255 ( .A1(n1359), .A2(n1361), .ZN(n3461) );
  NAND2_X1 U3256 ( .A1(n1384), .A2(n1361), .ZN(n3462) );
  NAND3_X1 U3257 ( .A1(n3460), .A2(n3462), .A3(n3461), .ZN(n1354) );
  NAND2_X1 U3258 ( .A1(n1559), .A2(n3464), .ZN(n3465) );
  NAND2_X1 U3259 ( .A1(n3463), .A2(n1557), .ZN(n3466) );
  NAND2_X1 U3260 ( .A1(n3465), .A2(n3466), .ZN(n3666) );
  INV_X1 U3261 ( .A(n1559), .ZN(n3463) );
  INV_X1 U3262 ( .A(n1557), .ZN(n3464) );
  NAND2_X1 U3263 ( .A1(n3716), .A2(n3468), .ZN(n3469) );
  NAND2_X1 U3264 ( .A1(n3467), .A2(n342), .ZN(n3470) );
  NAND2_X1 U3265 ( .A1(n3469), .A2(n3470), .ZN(n3236) );
  INV_X1 U3266 ( .A(n3716), .ZN(n3467) );
  INV_X1 U3267 ( .A(n342), .ZN(n3468) );
  INV_X1 U3268 ( .A(n712), .ZN(n710) );
  OAI21_X2 U3269 ( .B1(n692), .B2(n712), .A(n693), .ZN(n691) );
  AOI21_X2 U3270 ( .B1(n995), .B2(n721), .A(n714), .ZN(n712) );
  INV_X1 U3271 ( .A(n716), .ZN(n714) );
  NAND2_X1 U3272 ( .A1(n995), .A2(n716), .ZN(n549) );
  NAND2_X2 U3273 ( .A1(n3232), .A2(n402), .ZN(n3509) );
  AND2_X2 U3274 ( .A1(n3236), .A2(n390), .ZN(n3725) );
  XNOR2_X1 U3275 ( .A(n1520), .B(n1493), .ZN(n3698) );
  NAND2_X2 U3276 ( .A1(n3489), .A2(n3490), .ZN(n2256) );
  AND2_X1 U3277 ( .A1(n3228), .A2(n3642), .ZN(n3690) );
  INV_X1 U3278 ( .A(n3799), .ZN(n3471) );
  AND2_X1 U3279 ( .A1(n3232), .A2(n402), .ZN(n3799) );
  AND2_X1 U3280 ( .A1(n3688), .A2(n3689), .ZN(n3472) );
  INV_X1 U3281 ( .A(n3795), .ZN(n3473) );
  INV_X1 U3282 ( .A(n3657), .ZN(n3474) );
  INV_X4 U3283 ( .A(a[4]), .ZN(n3583) );
  INV_X4 U3284 ( .A(n3798), .ZN(n3721) );
  NOR2_X1 U3285 ( .A1(n1820), .A2(n1841), .ZN(n861) );
  INV_X1 U3286 ( .A(n3776), .ZN(n399) );
  NOR2_X2 U3287 ( .A1(n1111), .A2(n1122), .ZN(n663) );
  NOR2_X2 U3288 ( .A1(n663), .A2(n660), .ZN(n658) );
  NAND2_X2 U3289 ( .A1(n658), .A2(n989), .ZN(n656) );
  AOI21_X2 U3290 ( .B1(n658), .B2(n667), .A(n659), .ZN(n657) );
  INV_X2 U3291 ( .A(n3734), .ZN(n3737) );
  XOR2_X1 U3292 ( .A(n1501), .B(n1503), .Z(n3476) );
  XOR2_X1 U3293 ( .A(n1528), .B(n3476), .Z(n1495) );
  NAND2_X1 U3294 ( .A1(n1528), .A2(n1501), .ZN(n3477) );
  NAND2_X1 U3295 ( .A1(n1528), .A2(n1503), .ZN(n3478) );
  NAND2_X1 U3296 ( .A1(n1501), .A2(n1503), .ZN(n3479) );
  NAND3_X1 U3297 ( .A1(n3477), .A2(n3479), .A3(n3478), .ZN(n1494) );
  NOR2_X1 U3298 ( .A1(n1698), .A2(n1723), .ZN(n824) );
  NAND2_X1 U3299 ( .A1(n1698), .A2(n1723), .ZN(n825) );
  OAI22_X1 U3300 ( .A1(n3709), .A2(n2907), .B1(n2906), .B2(n393), .ZN(n2341)
         );
  OAI22_X1 U3301 ( .A1(n3708), .A2(n3284), .B1(n2931), .B2(n393), .ZN(n2068)
         );
  OAI22_X1 U3302 ( .A1(n3709), .A2(n2906), .B1(n2905), .B2(n393), .ZN(n2340)
         );
  OAI22_X1 U3303 ( .A1(n3709), .A2(n2925), .B1(n2924), .B2(n393), .ZN(n2359)
         );
  OAI22_X1 U3304 ( .A1(n3708), .A2(n2899), .B1(n393), .B2(n3284), .ZN(n2333)
         );
  OAI22_X1 U3305 ( .A1(n3709), .A2(n2924), .B1(n2923), .B2(n393), .ZN(n2358)
         );
  OAI22_X1 U3306 ( .A1(n3708), .A2(n2920), .B1(n2919), .B2(n393), .ZN(n2354)
         );
  OAI22_X1 U3307 ( .A1(n443), .A2(n2914), .B1(n2913), .B2(n393), .ZN(n2348) );
  OAI22_X1 U3308 ( .A1(n3709), .A2(n2918), .B1(n2917), .B2(n393), .ZN(n2352)
         );
  OAI22_X1 U3309 ( .A1(n443), .A2(n2922), .B1(n2921), .B2(n393), .ZN(n2356) );
  NOR2_X1 U3310 ( .A1(n699), .A2(n696), .ZN(n3480) );
  NOR2_X2 U3311 ( .A1(n699), .A2(n696), .ZN(n694) );
  XOR2_X1 U3312 ( .A(n2544), .B(n2416), .Z(n3481) );
  XOR2_X1 U3313 ( .A(n3481), .B(n2256), .Z(n1690) );
  XOR2_X1 U3314 ( .A(n1692), .B(n1694), .Z(n3482) );
  XOR2_X1 U3315 ( .A(n3482), .B(n1690), .Z(n1680) );
  NAND2_X1 U3316 ( .A1(n2544), .A2(n2416), .ZN(n3483) );
  NAND2_X1 U3317 ( .A1(n2544), .A2(n2256), .ZN(n3484) );
  NAND2_X1 U3318 ( .A1(n2416), .A2(n2256), .ZN(n3485) );
  NAND3_X1 U3319 ( .A1(n3483), .A2(n3484), .A3(n3485), .ZN(n1689) );
  NAND2_X1 U3320 ( .A1(n1692), .A2(n1694), .ZN(n3486) );
  NAND2_X1 U3321 ( .A1(n1692), .A2(n1690), .ZN(n3487) );
  NAND2_X1 U3322 ( .A1(n1694), .A2(n1690), .ZN(n3488) );
  NAND3_X1 U3323 ( .A1(n3486), .A2(n3487), .A3(n3488), .ZN(n1679) );
  OR2_X1 U3324 ( .A1(n3779), .A2(n2825), .ZN(n3489) );
  OR2_X1 U3325 ( .A1(n2824), .A2(n402), .ZN(n3490) );
  XNOR2_X1 U3326 ( .A(n479), .B(n354), .ZN(n2825) );
  XNOR2_X1 U3327 ( .A(n481), .B(n354), .ZN(n2824) );
  INV_X1 U3328 ( .A(n696), .ZN(n992) );
  OAI21_X1 U3329 ( .B1(n696), .B2(n700), .A(n697), .ZN(n695) );
  NAND2_X1 U3330 ( .A1(n1167), .A2(n1182), .ZN(n697) );
  INV_X8 U3331 ( .A(n3803), .ZN(n3491) );
  OR2_X1 U3332 ( .A1(n446), .A2(n2879), .ZN(n3492) );
  OR2_X1 U3333 ( .A1(n2878), .A2(n3729), .ZN(n3493) );
  NAND2_X1 U3334 ( .A1(n3492), .A2(n3493), .ZN(n2312) );
  INV_X4 U3335 ( .A(n3803), .ZN(n446) );
  XNOR2_X1 U3336 ( .A(n503), .B(n348), .ZN(n2879) );
  XNOR2_X1 U3337 ( .A(n505), .B(n348), .ZN(n2878) );
  INV_X4 U3338 ( .A(n3732), .ZN(n3494) );
  INV_X4 U3339 ( .A(n3732), .ZN(n434) );
  NAND2_X1 U3340 ( .A1(n635), .A2(n676), .ZN(n3495) );
  INV_X1 U3341 ( .A(n636), .ZN(n3496) );
  AND2_X2 U3342 ( .A1(n3495), .A2(n3496), .ZN(n634) );
  OAI21_X1 U3343 ( .B1(n677), .B2(n681), .A(n678), .ZN(n676) );
  OAI21_X2 U3344 ( .B1(n634), .B2(n617), .A(n618), .ZN(n616) );
  BUF_X1 U3345 ( .A(n772), .Z(n3497) );
  INV_X4 U3346 ( .A(a[18]), .ZN(n3606) );
  INV_X2 U3347 ( .A(n3810), .ZN(n431) );
  AND2_X2 U3348 ( .A1(n3239), .A2(n3655), .ZN(n3810) );
  NAND2_X2 U3349 ( .A1(n1882), .A2(n1899), .ZN(n875) );
  NOR2_X1 U3350 ( .A1(n1882), .A2(n1899), .ZN(n874) );
  OAI22_X1 U3351 ( .A1(n443), .A2(n2929), .B1(n2928), .B2(n393), .ZN(n2363) );
  NAND2_X2 U3352 ( .A1(n3235), .A2(n393), .ZN(n3709) );
  OAI22_X1 U3353 ( .A1(n3709), .A2(n2926), .B1(n2925), .B2(n393), .ZN(n2360)
         );
  OAI22_X1 U3354 ( .A1(n3708), .A2(n2915), .B1(n2914), .B2(n393), .ZN(n2349)
         );
  OAI22_X1 U3355 ( .A1(n3708), .A2(n2916), .B1(n2915), .B2(n393), .ZN(n2350)
         );
  OAI22_X1 U3356 ( .A1(n3708), .A2(n2901), .B1(n2900), .B2(n393), .ZN(n2335)
         );
  OAI22_X1 U3357 ( .A1(n3709), .A2(n2905), .B1(n2904), .B2(n393), .ZN(n2339)
         );
  OAI22_X1 U3358 ( .A1(n3708), .A2(n2930), .B1(n2929), .B2(n393), .ZN(n2364)
         );
  OAI22_X1 U3359 ( .A1(n3708), .A2(n2927), .B1(n2926), .B2(n393), .ZN(n2361)
         );
  OAI22_X1 U3360 ( .A1(n443), .A2(n2921), .B1(n2920), .B2(n393), .ZN(n2355) );
  OAI22_X1 U3361 ( .A1(n3590), .A2(n3190), .B1(n3189), .B2(n369), .ZN(n2632)
         );
  OAI22_X1 U3362 ( .A1(n3590), .A2(n3186), .B1(n3185), .B2(n369), .ZN(n2628)
         );
  OAI22_X1 U3363 ( .A1(n3590), .A2(n3193), .B1(n3192), .B2(n369), .ZN(n2635)
         );
  OAI22_X1 U3364 ( .A1(n3590), .A2(n3194), .B1(n3193), .B2(n369), .ZN(n2636)
         );
  OAI22_X1 U3365 ( .A1(n3590), .A2(n3292), .B1(n3195), .B2(n369), .ZN(n2076)
         );
  OAI22_X1 U3366 ( .A1(n3590), .A2(n3191), .B1(n3190), .B2(n369), .ZN(n2633)
         );
  OAI22_X1 U3367 ( .A1(n3590), .A2(n3192), .B1(n3191), .B2(n369), .ZN(n2634)
         );
  OAI22_X1 U3368 ( .A1(n3590), .A2(n3189), .B1(n3188), .B2(n369), .ZN(n2631)
         );
  OAI22_X1 U3369 ( .A1(n3590), .A2(n3188), .B1(n3187), .B2(n369), .ZN(n2630)
         );
  OAI22_X1 U3370 ( .A1(n3590), .A2(n3187), .B1(n3186), .B2(n369), .ZN(n2629)
         );
  OAI22_X1 U3371 ( .A1(n3590), .A2(n3185), .B1(n3184), .B2(n369), .ZN(n2627)
         );
  OAI22_X1 U3372 ( .A1(n3590), .A2(n3178), .B1(n3177), .B2(n369), .ZN(n2620)
         );
  OAI22_X1 U3373 ( .A1(n3590), .A2(n3184), .B1(n3183), .B2(n369), .ZN(n2626)
         );
  OAI22_X1 U3374 ( .A1(n3590), .A2(n3183), .B1(n3182), .B2(n369), .ZN(n2625)
         );
  OAI22_X1 U3375 ( .A1(n3590), .A2(n3179), .B1(n3178), .B2(n369), .ZN(n2621)
         );
  OAI22_X1 U3376 ( .A1(n3590), .A2(n3164), .B1(n3163), .B2(n369), .ZN(n2606)
         );
  OAI22_X1 U3377 ( .A1(n3590), .A2(n3163), .B1(n3292), .B2(n369), .ZN(n2605)
         );
  OAI22_X1 U3378 ( .A1(n3590), .A2(n3181), .B1(n3180), .B2(n369), .ZN(n2623)
         );
  OAI22_X1 U3379 ( .A1(n3590), .A2(n3182), .B1(n3181), .B2(n369), .ZN(n2624)
         );
  OAI22_X1 U3380 ( .A1(n3590), .A2(n3176), .B1(n3175), .B2(n369), .ZN(n2618)
         );
  OAI22_X1 U3381 ( .A1(n3590), .A2(n3168), .B1(n3167), .B2(n369), .ZN(n2610)
         );
  OAI22_X1 U3382 ( .A1(n3598), .A2(n2975), .B1(n2974), .B2(n3736), .ZN(n2411)
         );
  OAI22_X1 U3383 ( .A1(n3598), .A2(n2969), .B1(n2968), .B2(n3737), .ZN(n2405)
         );
  OAI22_X1 U3384 ( .A1(n3598), .A2(n2992), .B1(n2991), .B2(n3737), .ZN(n2428)
         );
  OAI22_X1 U3385 ( .A1(n3598), .A2(n2968), .B1(n2967), .B2(n3737), .ZN(n2404)
         );
  OAI22_X1 U3386 ( .A1(n3598), .A2(n2965), .B1(n3736), .B2(n3286), .ZN(n2401)
         );
  OAI22_X1 U3387 ( .A1(n3598), .A2(n2977), .B1(n2976), .B2(n3737), .ZN(n2413)
         );
  OAI22_X1 U3388 ( .A1(n3598), .A2(n2966), .B1(n2965), .B2(n3736), .ZN(n2402)
         );
  OAI22_X1 U3389 ( .A1(n3598), .A2(n2967), .B1(n2966), .B2(n3736), .ZN(n2403)
         );
  OAI22_X1 U3390 ( .A1(n3598), .A2(n2987), .B1(n2986), .B2(n3736), .ZN(n2423)
         );
  OAI22_X1 U3391 ( .A1(n3598), .A2(n2996), .B1(n2995), .B2(n3736), .ZN(n2432)
         );
  OAI22_X1 U3392 ( .A1(n3598), .A2(n2991), .B1(n2990), .B2(n3736), .ZN(n2427)
         );
  OAI22_X1 U3393 ( .A1(n3598), .A2(n2990), .B1(n2989), .B2(n3737), .ZN(n2426)
         );
  OAI22_X1 U3394 ( .A1(n3598), .A2(n3286), .B1(n2997), .B2(n3737), .ZN(n2070)
         );
  OAI22_X1 U3395 ( .A1(n3598), .A2(n2995), .B1(n2994), .B2(n3736), .ZN(n2431)
         );
  OAI22_X1 U3396 ( .A1(n3598), .A2(n2994), .B1(n2993), .B2(n3737), .ZN(n2430)
         );
  INV_X2 U3397 ( .A(n3734), .ZN(n3736) );
  NAND2_X2 U3398 ( .A1(n3235), .A2(n393), .ZN(n443) );
  XNOR2_X1 U3399 ( .A(n3498), .B(n2218), .ZN(n1513) );
  XNOR2_X1 U3400 ( .A(n2186), .B(n2410), .ZN(n3498) );
  XOR2_X2 U3401 ( .A(n3499), .B(n1406), .Z(n1379) );
  NOR2_X2 U3402 ( .A1(n1183), .A2(n1200), .ZN(n699) );
  XOR2_X1 U3403 ( .A(n1383), .B(n1408), .Z(n3499) );
  XOR2_X1 U3404 ( .A(n1404), .B(n1381), .Z(n3500) );
  XOR2_X1 U3405 ( .A(n3500), .B(n1379), .Z(n1377) );
  NAND2_X1 U3406 ( .A1(n1383), .A2(n1408), .ZN(n3501) );
  NAND2_X1 U3407 ( .A1(n1383), .A2(n1406), .ZN(n3502) );
  NAND2_X1 U3408 ( .A1(n1408), .A2(n1406), .ZN(n3503) );
  NAND3_X1 U3409 ( .A1(n3501), .A2(n3502), .A3(n3503), .ZN(n1378) );
  NAND2_X1 U3410 ( .A1(n1404), .A2(n1381), .ZN(n3504) );
  NAND2_X1 U3411 ( .A1(n1404), .A2(n1379), .ZN(n3505) );
  NAND2_X1 U3412 ( .A1(n1381), .A2(n1379), .ZN(n3506) );
  NAND3_X1 U3413 ( .A1(n3504), .A2(n3505), .A3(n3506), .ZN(n1376) );
  XOR2_X1 U3414 ( .A(a[18]), .B(n348), .Z(n3234) );
  OAI22_X1 U3415 ( .A1(n3619), .A2(n3084), .B1(n3083), .B2(n3679), .ZN(n2523)
         );
  OAI22_X1 U3416 ( .A1(n3619), .A2(n3086), .B1(n3085), .B2(n3679), .ZN(n2525)
         );
  OAI22_X1 U3417 ( .A1(n3619), .A2(n3078), .B1(n3077), .B2(n3679), .ZN(n2517)
         );
  OAI22_X1 U3418 ( .A1(n3619), .A2(n3083), .B1(n3082), .B2(n3679), .ZN(n2522)
         );
  OAI22_X1 U3419 ( .A1(n3619), .A2(n3081), .B1(n3080), .B2(n3679), .ZN(n2520)
         );
  OAI22_X1 U3420 ( .A1(n3598), .A2(n2971), .B1(n2970), .B2(n3737), .ZN(n2407)
         );
  AND2_X2 U3421 ( .A1(n3232), .A2(n402), .ZN(n3507) );
  NAND2_X1 U3422 ( .A1(n3232), .A2(n402), .ZN(n3508) );
  XOR2_X1 U3423 ( .A(n1671), .B(n1646), .Z(n3510) );
  XOR2_X1 U3424 ( .A(n1644), .B(n3510), .Z(n1642) );
  NAND2_X1 U3425 ( .A1(n1644), .A2(n1671), .ZN(n3511) );
  NAND2_X1 U3426 ( .A1(n1644), .A2(n1646), .ZN(n3512) );
  NAND2_X1 U3427 ( .A1(n1671), .A2(n1646), .ZN(n3513) );
  NAND3_X1 U3428 ( .A1(n3511), .A2(n3513), .A3(n3512), .ZN(n1641) );
  XOR2_X2 U3429 ( .A(n3540), .B(n354), .Z(n3232) );
  BUF_X1 U3430 ( .A(n3604), .Z(n3514) );
  BUF_X1 U3431 ( .A(n997), .Z(n3515) );
  AND2_X2 U3432 ( .A1(n1281), .A2(n1302), .ZN(n3665) );
  NOR2_X1 U3433 ( .A1(n1259), .A2(n1280), .ZN(n735) );
  OAI22_X1 U3434 ( .A1(n3619), .A2(n3073), .B1(n3072), .B2(n3679), .ZN(n2512)
         );
  XOR2_X1 U3435 ( .A(n2385), .B(n2449), .Z(n3516) );
  XOR2_X1 U3436 ( .A(n3516), .B(n2417), .Z(n1714) );
  XOR2_X1 U3437 ( .A(n1741), .B(n1739), .Z(n3517) );
  XOR2_X1 U3438 ( .A(n3517), .B(n1714), .Z(n1710) );
  NAND2_X1 U3439 ( .A1(n2385), .A2(n2449), .ZN(n3518) );
  NAND2_X1 U3440 ( .A1(n2385), .A2(n2417), .ZN(n3519) );
  NAND2_X1 U3441 ( .A1(n2449), .A2(n2417), .ZN(n3520) );
  NAND3_X1 U3442 ( .A1(n3518), .A2(n3519), .A3(n3520), .ZN(n1713) );
  NAND2_X1 U3443 ( .A1(n1741), .A2(n1739), .ZN(n3521) );
  NAND2_X1 U3444 ( .A1(n1741), .A2(n1714), .ZN(n3522) );
  NAND2_X1 U3445 ( .A1(n1739), .A2(n1714), .ZN(n3523) );
  NAND3_X1 U3446 ( .A1(n3521), .A2(n3522), .A3(n3523), .ZN(n1709) );
  OR2_X1 U3447 ( .A1(n3598), .A2(n2981), .ZN(n3524) );
  OR2_X1 U3448 ( .A1(n2980), .A2(n3736), .ZN(n3525) );
  NAND2_X1 U3449 ( .A1(n3524), .A2(n3525), .ZN(n2417) );
  XNOR2_X1 U3450 ( .A(n497), .B(n339), .ZN(n2981) );
  XNOR2_X1 U3451 ( .A(n499), .B(n339), .ZN(n2980) );
  NOR2_X2 U3452 ( .A1(n788), .A2(n3754), .ZN(n786) );
  INV_X1 U3453 ( .A(n3665), .ZN(n739) );
  INV_X1 U3454 ( .A(n3643), .ZN(n738) );
  OAI21_X2 U3455 ( .B1(n877), .B2(n857), .A(n858), .ZN(n856) );
  XOR2_X1 U3456 ( .A(n2444), .B(n2220), .Z(n3526) );
  XOR2_X1 U3457 ( .A(n2252), .B(n3526), .Z(n1575) );
  NAND2_X1 U3458 ( .A1(n2252), .A2(n2444), .ZN(n3527) );
  NAND2_X1 U3459 ( .A1(n2252), .A2(n2220), .ZN(n3528) );
  NAND2_X1 U3460 ( .A1(n2444), .A2(n2220), .ZN(n3529) );
  NAND3_X1 U3461 ( .A1(n3527), .A2(n3529), .A3(n3528), .ZN(n1574) );
  OR2_X1 U3462 ( .A1(n3509), .A2(n2821), .ZN(n3530) );
  OR2_X1 U3463 ( .A1(n2820), .A2(n402), .ZN(n3531) );
  NAND2_X1 U3464 ( .A1(n3530), .A2(n3531), .ZN(n2252) );
  OAI22_X1 U3465 ( .A1(n3706), .A2(n2790), .B1(n2789), .B2(n3581), .ZN(n2220)
         );
  XNOR2_X1 U3466 ( .A(n487), .B(n354), .ZN(n2821) );
  XNOR2_X1 U3467 ( .A(n489), .B(n354), .ZN(n2820) );
  INV_X1 U3468 ( .A(n735), .ZN(n997) );
  XNOR2_X2 U3469 ( .A(n3724), .B(n3278), .ZN(n3532) );
  INV_X4 U3470 ( .A(n3532), .ZN(n3791) );
  INV_X4 U3471 ( .A(n363), .ZN(n3278) );
  XOR2_X1 U3472 ( .A(n1509), .B(n1517), .Z(n3533) );
  XOR2_X1 U3473 ( .A(n1540), .B(n3533), .Z(n1503) );
  NAND2_X1 U3474 ( .A1(n1540), .A2(n1509), .ZN(n3534) );
  NAND2_X1 U3475 ( .A1(n1540), .A2(n1517), .ZN(n3535) );
  NAND2_X1 U3476 ( .A1(n1509), .A2(n1517), .ZN(n3536) );
  NAND3_X1 U3477 ( .A1(n3534), .A2(n3536), .A3(n3535), .ZN(n1502) );
  BUF_X1 U3478 ( .A(n3756), .Z(n3537) );
  NOR2_X1 U3479 ( .A1(n1431), .A2(n1458), .ZN(n3756) );
  NAND2_X2 U3480 ( .A1(n3235), .A2(n393), .ZN(n3708) );
  OAI22_X1 U3481 ( .A1(n443), .A2(n2909), .B1(n2908), .B2(n393), .ZN(n2343) );
  OAI22_X1 U3482 ( .A1(n3708), .A2(n2928), .B1(n2927), .B2(n393), .ZN(n2362)
         );
  OAI22_X1 U3483 ( .A1(n3708), .A2(n2902), .B1(n2901), .B2(n393), .ZN(n2336)
         );
  OAI22_X1 U3484 ( .A1(n3709), .A2(n2900), .B1(n2899), .B2(n393), .ZN(n2334)
         );
  OAI22_X1 U3485 ( .A1(n3709), .A2(n2903), .B1(n2902), .B2(n393), .ZN(n2337)
         );
  OAI22_X1 U3486 ( .A1(n3709), .A2(n2904), .B1(n2903), .B2(n393), .ZN(n2338)
         );
  OAI22_X1 U3487 ( .A1(n3708), .A2(n2917), .B1(n2916), .B2(n393), .ZN(n2351)
         );
  OAI22_X1 U3488 ( .A1(n3709), .A2(n2919), .B1(n2918), .B2(n393), .ZN(n2353)
         );
  OAI22_X1 U3489 ( .A1(n3709), .A2(n2923), .B1(n2922), .B2(n393), .ZN(n2357)
         );
  OAI22_X1 U3490 ( .A1(n3708), .A2(n2912), .B1(n2911), .B2(n393), .ZN(n2346)
         );
  XNOR2_X1 U3491 ( .A(n3538), .B(n1794), .ZN(n1782) );
  XNOR2_X1 U3492 ( .A(n1790), .B(n1792), .ZN(n3538) );
  OAI22_X1 U3493 ( .A1(n446), .A2(n2877), .B1(n2876), .B2(n3729), .ZN(n2310)
         );
  XNOR2_X2 U3494 ( .A(a[8]), .B(n3289), .ZN(n3539) );
  INV_X2 U3495 ( .A(n3588), .ZN(n3798) );
  OAI22_X1 U3496 ( .A1(n437), .A2(n2984), .B1(n2983), .B2(n3736), .ZN(n2420)
         );
  OAI22_X1 U3497 ( .A1(n437), .A2(n2986), .B1(n2985), .B2(n3737), .ZN(n2422)
         );
  OAI22_X1 U3498 ( .A1(n437), .A2(n2989), .B1(n2988), .B2(n3737), .ZN(n2425)
         );
  OAI22_X1 U3499 ( .A1(n437), .A2(n2985), .B1(n2984), .B2(n3736), .ZN(n2421)
         );
  OAI22_X1 U3500 ( .A1(n437), .A2(n2973), .B1(n2972), .B2(n3737), .ZN(n2409)
         );
  OAI22_X1 U3501 ( .A1(n437), .A2(n2980), .B1(n2979), .B2(n3736), .ZN(n2416)
         );
  OAI22_X1 U3502 ( .A1(n437), .A2(n2970), .B1(n2969), .B2(n3737), .ZN(n2406)
         );
  OAI22_X1 U3503 ( .A1(n437), .A2(n2979), .B1(n2978), .B2(n3736), .ZN(n2415)
         );
  BUF_X1 U3504 ( .A(a[22]), .Z(n3540) );
  XOR2_X1 U3505 ( .A(n1378), .B(n1355), .Z(n3541) );
  XOR2_X2 U3506 ( .A(n1353), .B(n3541), .Z(n1351) );
  NAND2_X1 U3507 ( .A1(n1353), .A2(n1378), .ZN(n3542) );
  NAND2_X1 U3508 ( .A1(n1353), .A2(n1355), .ZN(n3543) );
  NAND2_X1 U3509 ( .A1(n1378), .A2(n1355), .ZN(n3544) );
  NAND3_X1 U3510 ( .A1(n3542), .A2(n3544), .A3(n3543), .ZN(n1350) );
  INV_X1 U3511 ( .A(n690), .ZN(n688) );
  OAI22_X1 U3512 ( .A1(n3598), .A2(n2993), .B1(n2992), .B2(n3736), .ZN(n2429)
         );
  NOR2_X2 U3513 ( .A1(n1934), .A2(n1949), .ZN(n890) );
  NAND2_X2 U3514 ( .A1(n1934), .A2(n1949), .ZN(n891) );
  XNOR2_X2 U3515 ( .A(n3572), .B(n324), .ZN(n3242) );
  INV_X4 U3516 ( .A(n3810), .ZN(n3793) );
  INV_X4 U3517 ( .A(n3777), .ZN(n3545) );
  AND2_X2 U3518 ( .A1(n3701), .A2(n3702), .ZN(n3589) );
  OAI21_X1 U3519 ( .B1(n805), .B2(n784), .A(n785), .ZN(n783) );
  NAND2_X1 U3520 ( .A1(n996), .A2(n995), .ZN(n711) );
  NAND2_X1 U3521 ( .A1(n996), .A2(n719), .ZN(n550) );
  INV_X1 U3522 ( .A(n718), .ZN(n996) );
  NOR2_X1 U3523 ( .A1(n1239), .A2(n1258), .ZN(n718) );
  NAND2_X2 U3524 ( .A1(n1239), .A2(n1258), .ZN(n719) );
  INV_X4 U3525 ( .A(n345), .ZN(n3546) );
  INV_X4 U3526 ( .A(n3546), .ZN(n3547) );
  NOR2_X2 U3527 ( .A1(n3654), .A2(n747), .ZN(n729) );
  OAI22_X1 U3528 ( .A1(n458), .A2(n2746), .B1(n2745), .B2(n3742), .ZN(n2175)
         );
  OAI22_X1 U3529 ( .A1(n458), .A2(n2761), .B1(n2760), .B2(n3742), .ZN(n2190)
         );
  OAI22_X1 U3530 ( .A1(n458), .A2(n2748), .B1(n2747), .B2(n3742), .ZN(n2177)
         );
  OAI22_X1 U3531 ( .A1(n458), .A2(n2765), .B1(n2764), .B2(n3741), .ZN(n2194)
         );
  OAI22_X1 U3532 ( .A1(n458), .A2(n2764), .B1(n2763), .B2(n3742), .ZN(n2193)
         );
  OAI22_X1 U3533 ( .A1(n458), .A2(n2760), .B1(n2759), .B2(n3741), .ZN(n2189)
         );
  OAI22_X1 U3534 ( .A1(n458), .A2(n2753), .B1(n2752), .B2(n3741), .ZN(n2182)
         );
  OAI22_X1 U3535 ( .A1(n458), .A2(n2755), .B1(n2754), .B2(n3741), .ZN(n2184)
         );
  OAI22_X1 U3536 ( .A1(n458), .A2(n2759), .B1(n2758), .B2(n3741), .ZN(n2188)
         );
  OAI22_X1 U3537 ( .A1(n458), .A2(n2754), .B1(n2753), .B2(n3741), .ZN(n2183)
         );
  OAI22_X1 U3538 ( .A1(n458), .A2(n2756), .B1(n2755), .B2(n3742), .ZN(n2185)
         );
  OAI22_X1 U3539 ( .A1(n458), .A2(n2762), .B1(n2761), .B2(n3741), .ZN(n2191)
         );
  NAND2_X1 U3540 ( .A1(n1303), .A2(n1326), .ZN(n748) );
  NOR2_X2 U3541 ( .A1(n1303), .A2(n1326), .ZN(n747) );
  INV_X1 U3542 ( .A(n345), .ZN(n3570) );
  BUF_X1 U3543 ( .A(n856), .Z(n3548) );
  INV_X4 U3544 ( .A(n3448), .ZN(n3549) );
  INV_X2 U3545 ( .A(n3549), .ZN(n3550) );
  XOR2_X1 U3546 ( .A(n2612), .B(n2420), .Z(n3551) );
  XOR2_X1 U3547 ( .A(n3551), .B(n2260), .Z(n1794) );
  NAND2_X1 U3548 ( .A1(n2612), .A2(n2420), .ZN(n3552) );
  NAND2_X1 U3549 ( .A1(n2612), .A2(n2260), .ZN(n3553) );
  NAND2_X1 U3550 ( .A1(n2420), .A2(n2260), .ZN(n3554) );
  NAND3_X1 U3551 ( .A1(n3552), .A2(n3553), .A3(n3554), .ZN(n1793) );
  NAND2_X1 U3552 ( .A1(n1790), .A2(n1792), .ZN(n3555) );
  NAND2_X1 U3553 ( .A1(n1790), .A2(n1794), .ZN(n3556) );
  NAND2_X1 U3554 ( .A1(n1792), .A2(n1794), .ZN(n3557) );
  NAND3_X1 U3555 ( .A1(n3555), .A2(n3556), .A3(n3557), .ZN(n1781) );
  OR2_X1 U3556 ( .A1(n2829), .A2(n3509), .ZN(n3558) );
  OR2_X1 U3557 ( .A1(n2828), .A2(n402), .ZN(n3559) );
  NAND2_X1 U3558 ( .A1(n3558), .A2(n3559), .ZN(n2260) );
  XNOR2_X1 U3559 ( .A(n471), .B(n354), .ZN(n2829) );
  XNOR2_X1 U3560 ( .A(n473), .B(n354), .ZN(n2828) );
  BUF_X1 U3561 ( .A(n815), .Z(n3560) );
  INV_X4 U3562 ( .A(n3806), .ZN(n3562) );
  INV_X4 U3563 ( .A(n3806), .ZN(n3561) );
  INV_X2 U3564 ( .A(n348), .ZN(n3563) );
  INV_X1 U3565 ( .A(n3806), .ZN(n449) );
  INV_X1 U3566 ( .A(n348), .ZN(n3283) );
  AND2_X4 U3567 ( .A1(n3233), .A2(n3612), .ZN(n3806) );
  OAI22_X1 U3568 ( .A1(n437), .A2(n2982), .B1(n2981), .B2(n3737), .ZN(n2418)
         );
  OAI21_X1 U3569 ( .B1(n819), .B2(n825), .A(n820), .ZN(n3564) );
  OAI21_X1 U3570 ( .B1(n819), .B2(n825), .A(n820), .ZN(n818) );
  BUF_X1 U3571 ( .A(n3509), .Z(n3565) );
  NAND2_X1 U3572 ( .A1(n851), .A2(n850), .ZN(n571) );
  INV_X1 U3573 ( .A(n850), .ZN(n852) );
  OAI21_X1 U3574 ( .B1(n855), .B2(n849), .A(n850), .ZN(n848) );
  NAND2_X1 U3575 ( .A1(n1798), .A2(n1819), .ZN(n850) );
  OAI22_X1 U3576 ( .A1(n3619), .A2(n3091), .B1(n3090), .B2(n3678), .ZN(n2530)
         );
  OAI22_X1 U3577 ( .A1(n3620), .A2(n3069), .B1(n3068), .B2(n3678), .ZN(n2508)
         );
  OAI22_X1 U3578 ( .A1(n3619), .A2(n3075), .B1(n3074), .B2(n3678), .ZN(n2514)
         );
  OAI22_X1 U3579 ( .A1(n3619), .A2(n3090), .B1(n3089), .B2(n3678), .ZN(n2529)
         );
  OAI22_X1 U3580 ( .A1(n3620), .A2(n3085), .B1(n3084), .B2(n3678), .ZN(n2524)
         );
  OAI22_X1 U3581 ( .A1(n3619), .A2(n3068), .B1(n3067), .B2(n3678), .ZN(n2507)
         );
  OAI22_X1 U3582 ( .A1(n3619), .A2(n3092), .B1(n3091), .B2(n3678), .ZN(n2531)
         );
  OAI22_X1 U3583 ( .A1(n3620), .A2(n3071), .B1(n3070), .B2(n3678), .ZN(n2510)
         );
  OAI22_X1 U3584 ( .A1(n3620), .A2(n3082), .B1(n3081), .B2(n3678), .ZN(n2521)
         );
  OAI22_X1 U3585 ( .A1(n3619), .A2(n3095), .B1(n3094), .B2(n3678), .ZN(n2534)
         );
  OAI22_X1 U3586 ( .A1(n3620), .A2(n3074), .B1(n3073), .B2(n3678), .ZN(n2513)
         );
  OAI22_X1 U3587 ( .A1(n3620), .A2(n3089), .B1(n3088), .B2(n3678), .ZN(n2528)
         );
  OAI22_X1 U3588 ( .A1(n3620), .A2(n3066), .B1(n3065), .B2(n3678), .ZN(n2505)
         );
  OAI22_X1 U3589 ( .A1(n3620), .A2(n3077), .B1(n3076), .B2(n3678), .ZN(n2516)
         );
  OAI22_X1 U3590 ( .A1(n428), .A2(n3076), .B1(n3075), .B2(n3678), .ZN(n2515)
         );
  XOR2_X1 U3591 ( .A(n1643), .B(n1616), .Z(n3566) );
  XOR2_X1 U3592 ( .A(n1614), .B(n3566), .Z(n1612) );
  NAND2_X1 U3593 ( .A1(n1614), .A2(n1643), .ZN(n3567) );
  NAND2_X1 U3594 ( .A1(n1614), .A2(n1616), .ZN(n3568) );
  NAND2_X1 U3595 ( .A1(n1643), .A2(n1616), .ZN(n3569) );
  NAND3_X1 U3596 ( .A1(n3567), .A2(n3569), .A3(n3568), .ZN(n1611) );
  OAI21_X4 U3597 ( .B1(n754), .B2(n760), .A(n755), .ZN(n753) );
  INV_X2 U3598 ( .A(n3570), .ZN(n3571) );
  INV_X8 U3599 ( .A(n3808), .ZN(n458) );
  INV_X8 U3600 ( .A(n3809), .ZN(n3573) );
  INV_X4 U3601 ( .A(n3809), .ZN(n372) );
  INV_X2 U3602 ( .A(n416), .ZN(n3574) );
  INV_X16 U3603 ( .A(n3574), .ZN(n3575) );
  INV_X4 U3604 ( .A(n366), .ZN(n416) );
  OR2_X2 U3605 ( .A1(n1750), .A2(n1773), .ZN(n3576) );
  NOR2_X1 U3606 ( .A1(n1950), .A2(n1963), .ZN(n902) );
  NAND2_X2 U3607 ( .A1(n1950), .A2(n1963), .ZN(n903) );
  AOI21_X2 U3608 ( .B1(n885), .B2(n893), .A(n886), .ZN(n884) );
  BUF_X1 U3609 ( .A(n804), .Z(n3577) );
  INV_X8 U3610 ( .A(n3725), .ZN(n3578) );
  INV_X4 U3611 ( .A(n3725), .ZN(n440) );
  AOI21_X2 U3612 ( .B1(n3438), .B2(n868), .A(n860), .ZN(n858) );
  OAI22_X1 U3613 ( .A1(n3598), .A2(n2988), .B1(n2987), .B2(n3736), .ZN(n2424)
         );
  NOR2_X1 U3614 ( .A1(n1612), .A2(n1641), .ZN(n3605) );
  NAND2_X1 U3615 ( .A1(n1010), .A2(n812), .ZN(n564) );
  INV_X2 U3616 ( .A(n3807), .ZN(n3796) );
  XNOR2_X2 U3617 ( .A(n1521), .B(n3675), .ZN(n1519) );
  INV_X4 U3618 ( .A(n3611), .ZN(n3613) );
  OAI22_X1 U3619 ( .A1(n3723), .A2(n3149), .B1(n3148), .B2(n3573), .ZN(n2590)
         );
  OAI22_X1 U3620 ( .A1(n3619), .A2(n3087), .B1(n3086), .B2(n3679), .ZN(n2526)
         );
  AND2_X1 U3621 ( .A1(n3231), .A2(n405), .ZN(n3579) );
  INV_X8 U3622 ( .A(n3800), .ZN(n3581) );
  INV_X1 U3623 ( .A(n3800), .ZN(n405) );
  NOR2_X2 U3624 ( .A1(n1842), .A2(n1861), .ZN(n864) );
  NAND2_X1 U3625 ( .A1(n1842), .A2(n1861), .ZN(n865) );
  INV_X1 U3626 ( .A(n803), .ZN(n1009) );
  INV_X1 U3627 ( .A(n798), .ZN(n796) );
  INV_X1 U3628 ( .A(n847), .ZN(n845) );
  NAND2_X1 U3629 ( .A1(n3773), .A2(n801), .ZN(n562) );
  NAND2_X1 U3630 ( .A1(n1551), .A2(n1581), .ZN(n801) );
  INV_X1 U3631 ( .A(n3589), .ZN(n3777) );
  NOR2_X1 U3632 ( .A1(n1431), .A2(n1458), .ZN(n777) );
  INV_X4 U3633 ( .A(n3810), .ZN(n3794) );
  INV_X2 U3634 ( .A(n806), .ZN(n805) );
  BUF_X1 U3635 ( .A(n706), .Z(n3582) );
  NAND2_X2 U3636 ( .A1(a[4]), .A2(n324), .ZN(n3585) );
  NAND2_X1 U3637 ( .A1(n3583), .A2(n3584), .ZN(n3586) );
  NAND2_X1 U3638 ( .A1(n3585), .A2(n3586), .ZN(n3684) );
  INV_X2 U3639 ( .A(n324), .ZN(n3584) );
  OAI21_X1 U3640 ( .B1(n604), .B2(n531), .A(n605), .ZN(n603) );
  OAI21_X1 U3641 ( .B1(n707), .B2(n531), .A(n708), .ZN(n706) );
  NAND2_X1 U3642 ( .A1(n1750), .A2(n1773), .ZN(n840) );
  INV_X4 U3643 ( .A(n3507), .ZN(n3778) );
  XNOR2_X2 U3644 ( .A(n3587), .B(n2440), .ZN(n1451) );
  XNOR2_X1 U3645 ( .A(n2408), .B(n2248), .ZN(n3587) );
  INV_X2 U3646 ( .A(n396), .ZN(n3726) );
  XNOR2_X2 U3647 ( .A(a[10]), .B(n333), .ZN(n3588) );
  AOI21_X1 U3648 ( .B1(n603), .B2(n980), .A(n600), .ZN(n598) );
  NAND2_X1 U3649 ( .A1(n611), .A2(n981), .ZN(n604) );
  NAND2_X1 U3650 ( .A1(n3643), .A2(n739), .ZN(n552) );
  INV_X1 U3651 ( .A(n727), .ZN(n725) );
  NOR2_X2 U3652 ( .A1(n727), .A2(n613), .ZN(n611) );
  NAND2_X1 U3653 ( .A1(n822), .A2(n825), .ZN(n567) );
  INV_X1 U3654 ( .A(n825), .ZN(n823) );
  OAI22_X1 U3655 ( .A1(n3704), .A2(n2798), .B1(n2797), .B2(n3581), .ZN(n2228)
         );
  NAND2_X4 U3656 ( .A1(n3243), .A2(n369), .ZN(n3590) );
  XNOR2_X1 U3657 ( .A(n529), .B(n321), .ZN(n3163) );
  XNOR2_X1 U3658 ( .A(n527), .B(n321), .ZN(n3164) );
  XNOR2_X1 U3659 ( .A(n525), .B(n321), .ZN(n3165) );
  XNOR2_X1 U3660 ( .A(n523), .B(n321), .ZN(n3166) );
  XNOR2_X1 U3661 ( .A(n521), .B(n321), .ZN(n3167) );
  XNOR2_X1 U3662 ( .A(n519), .B(n321), .ZN(n3168) );
  XNOR2_X1 U3663 ( .A(n517), .B(n321), .ZN(n3169) );
  XNOR2_X1 U3664 ( .A(n515), .B(n321), .ZN(n3170) );
  XNOR2_X1 U3665 ( .A(n513), .B(n321), .ZN(n3171) );
  XNOR2_X1 U3666 ( .A(n511), .B(n321), .ZN(n3172) );
  XNOR2_X1 U3667 ( .A(n509), .B(n321), .ZN(n3173) );
  XNOR2_X1 U3668 ( .A(n483), .B(n321), .ZN(n3186) );
  XNOR2_X1 U3669 ( .A(n481), .B(n321), .ZN(n3187) );
  XNOR2_X1 U3670 ( .A(n479), .B(n321), .ZN(n3188) );
  XNOR2_X1 U3671 ( .A(n485), .B(n321), .ZN(n3185) );
  XNOR2_X1 U3672 ( .A(n487), .B(n321), .ZN(n3184) );
  XNOR2_X1 U3673 ( .A(n489), .B(n321), .ZN(n3183) );
  XNOR2_X1 U3674 ( .A(n491), .B(n321), .ZN(n3182) );
  XNOR2_X1 U3675 ( .A(n493), .B(n321), .ZN(n3181) );
  XNOR2_X1 U3676 ( .A(n495), .B(n321), .ZN(n3180) );
  XNOR2_X1 U3677 ( .A(n497), .B(n321), .ZN(n3179) );
  XNOR2_X1 U3678 ( .A(n499), .B(n321), .ZN(n3178) );
  XNOR2_X1 U3679 ( .A(n501), .B(n321), .ZN(n3177) );
  XNOR2_X1 U3680 ( .A(n503), .B(n321), .ZN(n3176) );
  XNOR2_X1 U3681 ( .A(n505), .B(n321), .ZN(n3175) );
  XNOR2_X1 U3682 ( .A(n507), .B(n321), .ZN(n3174) );
  BUF_X1 U3683 ( .A(n321), .Z(n3640) );
  XNOR2_X1 U3684 ( .A(a[20]), .B(n3563), .ZN(n3776) );
  INV_X1 U3685 ( .A(n3590), .ZN(n3813) );
  XOR2_X1 U3686 ( .A(n1511), .B(n1515), .Z(n3591) );
  XOR2_X1 U3687 ( .A(n3591), .B(n1513), .Z(n1501) );
  NAND2_X1 U3688 ( .A1(n2186), .A2(n2410), .ZN(n3592) );
  NAND2_X2 U3689 ( .A1(n2186), .A2(n2218), .ZN(n3593) );
  NAND2_X1 U3690 ( .A1(n2410), .A2(n2218), .ZN(n3594) );
  NAND3_X1 U3691 ( .A1(n3592), .A2(n3593), .A3(n3594), .ZN(n1512) );
  NAND2_X1 U3692 ( .A1(n1511), .A2(n1515), .ZN(n3595) );
  NAND2_X1 U3693 ( .A1(n1511), .A2(n1513), .ZN(n3596) );
  NAND2_X1 U3694 ( .A1(n1515), .A2(n1513), .ZN(n3597) );
  NAND3_X1 U3695 ( .A1(n3595), .A2(n3596), .A3(n3597), .ZN(n1500) );
  INV_X8 U3696 ( .A(n3805), .ZN(n3598) );
  AND2_X4 U3697 ( .A1(n3237), .A2(n3735), .ZN(n3805) );
  INV_X4 U3698 ( .A(n3805), .ZN(n437) );
  NAND2_X2 U3699 ( .A1(n775), .A2(n767), .ZN(n765) );
  INV_X1 U3700 ( .A(n840), .ZN(n838) );
  NAND2_X1 U3701 ( .A1(n3599), .A2(n3600), .ZN(n3602) );
  NAND2_X1 U3702 ( .A1(n3601), .A2(n3602), .ZN(n3663) );
  INV_X2 U3703 ( .A(n342), .ZN(n3600) );
  INV_X2 U3704 ( .A(n3468), .ZN(n3603) );
  INV_X8 U3705 ( .A(n3747), .ZN(n402) );
  OR2_X2 U3706 ( .A1(n1724), .A2(n1749), .ZN(n3604) );
  NOR2_X1 U3707 ( .A1(n1377), .A2(n1402), .ZN(n3781) );
  NOR2_X1 U3708 ( .A1(n1377), .A2(n1402), .ZN(n769) );
  OAI22_X1 U3709 ( .A1(n3709), .A2(n2910), .B1(n2909), .B2(n393), .ZN(n2344)
         );
  NAND2_X1 U3710 ( .A1(n3607), .A2(a[18]), .ZN(n3608) );
  NAND2_X1 U3711 ( .A1(n3608), .A2(n3609), .ZN(n3789) );
  INV_X2 U3712 ( .A(n345), .ZN(n3607) );
  NOR2_X1 U3713 ( .A1(n1612), .A2(n1641), .ZN(n811) );
  XNOR2_X1 U3714 ( .A(n3610), .B(n2187), .ZN(n1543) );
  XNOR2_X1 U3715 ( .A(n3634), .B(n2507), .ZN(n3610) );
  OAI22_X1 U3716 ( .A1(n3491), .A2(n2888), .B1(n2887), .B2(n3729), .ZN(n2321)
         );
  AND2_X2 U3717 ( .A1(n3229), .A2(n3589), .ZN(n3807) );
  OAI22_X1 U3718 ( .A1(n3491), .A2(n2881), .B1(n2880), .B2(n3728), .ZN(n2314)
         );
  INV_X1 U3719 ( .A(n3703), .ZN(n375) );
  OAI22_X1 U3720 ( .A1(n3706), .A2(n2785), .B1(n2784), .B2(n3581), .ZN(n2215)
         );
  OAI22_X1 U3721 ( .A1(n3704), .A2(n2788), .B1(n2787), .B2(n3581), .ZN(n2218)
         );
  INV_X1 U3722 ( .A(n3611), .ZN(n3612) );
  NOR2_X1 U3723 ( .A1(n3721), .A2(n3444), .ZN(n2467) );
  OAI22_X1 U3724 ( .A1(n3494), .A2(n2999), .B1(n2998), .B2(n3721), .ZN(n2436)
         );
  OAI22_X1 U3725 ( .A1(n3494), .A2(n3016), .B1(n3015), .B2(n3721), .ZN(n2453)
         );
  OAI22_X1 U3726 ( .A1(n3494), .A2(n3029), .B1(n3028), .B2(n3721), .ZN(n2466)
         );
  OAI22_X1 U3727 ( .A1(n3494), .A2(n3011), .B1(n3010), .B2(n3721), .ZN(n2448)
         );
  OAI22_X1 U3728 ( .A1(n3494), .A2(n3287), .B1(n3030), .B2(n3721), .ZN(n2071)
         );
  OAI22_X1 U3729 ( .A1(n3494), .A2(n3000), .B1(n2999), .B2(n3721), .ZN(n2437)
         );
  OAI22_X1 U3730 ( .A1(n3494), .A2(n3010), .B1(n3009), .B2(n3721), .ZN(n2447)
         );
  OAI22_X1 U3731 ( .A1(n3494), .A2(n3023), .B1(n3022), .B2(n3721), .ZN(n2460)
         );
  OAI22_X1 U3732 ( .A1(n3494), .A2(n3008), .B1(n3007), .B2(n3721), .ZN(n2445)
         );
  OAI22_X1 U3733 ( .A1(n3494), .A2(n3028), .B1(n3027), .B2(n3721), .ZN(n2465)
         );
  OAI22_X1 U3734 ( .A1(n434), .A2(n3002), .B1(n3001), .B2(n3721), .ZN(n2439)
         );
  OAI22_X1 U3735 ( .A1(n3494), .A2(n3025), .B1(n3024), .B2(n3721), .ZN(n2462)
         );
  OAI22_X1 U3736 ( .A1(n3494), .A2(n3014), .B1(n3013), .B2(n3721), .ZN(n2451)
         );
  OAI22_X1 U3737 ( .A1(n3494), .A2(n3001), .B1(n3000), .B2(n3721), .ZN(n2438)
         );
  OAI22_X1 U3738 ( .A1(n3494), .A2(n3027), .B1(n3026), .B2(n3721), .ZN(n2464)
         );
  OAI22_X1 U3739 ( .A1(n3494), .A2(n3004), .B1(n3003), .B2(n3721), .ZN(n2441)
         );
  INV_X4 U3740 ( .A(n3808), .ZN(n3614) );
  NAND2_X1 U3741 ( .A1(a[26]), .A2(n3616), .ZN(n3617) );
  NAND2_X1 U3742 ( .A1(n3615), .A2(n357), .ZN(n3618) );
  INV_X2 U3743 ( .A(n357), .ZN(n3616) );
  INV_X1 U3744 ( .A(n3605), .ZN(n1010) );
  NOR2_X2 U3745 ( .A1(n1798), .A2(n1819), .ZN(n849) );
  INV_X8 U3746 ( .A(n3802), .ZN(n3620) );
  INV_X4 U3747 ( .A(n3802), .ZN(n3619) );
  INV_X1 U3748 ( .A(n3802), .ZN(n428) );
  AND2_X4 U3749 ( .A1(n3240), .A2(n3677), .ZN(n3802) );
  NOR2_X2 U3750 ( .A1(n814), .A2(n811), .ZN(n809) );
  NAND2_X1 U3751 ( .A1(n1583), .A2(n3622), .ZN(n3623) );
  NAND2_X1 U3752 ( .A1(n3621), .A2(n1555), .ZN(n3624) );
  NAND2_X1 U3753 ( .A1(n3623), .A2(n3624), .ZN(n3667) );
  INV_X1 U3754 ( .A(n1583), .ZN(n3621) );
  INV_X1 U3755 ( .A(n1555), .ZN(n3622) );
  INV_X4 U3756 ( .A(n3804), .ZN(n3626) );
  INV_X4 U3757 ( .A(n3804), .ZN(n3625) );
  INV_X1 U3758 ( .A(n3804), .ZN(n390) );
  XOR2_X1 U3759 ( .A(n1541), .B(n1545), .Z(n3627) );
  XOR2_X1 U3760 ( .A(n3627), .B(n1543), .Z(n1531) );
  NAND2_X1 U3761 ( .A1(n3634), .A2(n2507), .ZN(n3628) );
  NAND2_X1 U3762 ( .A1(n3634), .A2(n2187), .ZN(n3629) );
  NAND2_X1 U3763 ( .A1(n2507), .A2(n2187), .ZN(n3630) );
  NAND3_X1 U3764 ( .A1(n3628), .A2(n3629), .A3(n3630), .ZN(n1542) );
  NAND2_X1 U3765 ( .A1(n1541), .A2(n1545), .ZN(n3631) );
  NAND2_X1 U3766 ( .A1(n1541), .A2(n1543), .ZN(n3632) );
  NAND2_X1 U3767 ( .A1(n1545), .A2(n1543), .ZN(n3633) );
  NAND3_X1 U3768 ( .A1(n3631), .A2(n3632), .A3(n3633), .ZN(n1530) );
  BUF_X2 U3769 ( .A(n2219), .Z(n3634) );
  OAI22_X1 U3770 ( .A1(n3705), .A2(n2789), .B1(n2788), .B2(n3581), .ZN(n2219)
         );
  OAI21_X1 U3771 ( .B1(n800), .B2(n3577), .A(n801), .ZN(n3635) );
  OAI21_X1 U3772 ( .B1(n804), .B2(n800), .A(n801), .ZN(n799) );
  OAI22_X1 U3773 ( .A1(n458), .A2(n2757), .B1(n2756), .B2(n3742), .ZN(n2186)
         );
  NAND2_X1 U3774 ( .A1(n3636), .A2(n3637), .ZN(n3639) );
  NAND2_X2 U3775 ( .A1(n3638), .A2(n3639), .ZN(n3809) );
  INV_X1 U3776 ( .A(n3572), .ZN(n3636) );
  OAI22_X1 U3777 ( .A1(n458), .A2(n2758), .B1(n2757), .B2(n3742), .ZN(n2187)
         );
  INV_X1 U3778 ( .A(n3733), .ZN(n387) );
  INV_X2 U3779 ( .A(n3472), .ZN(n3733) );
  OAI22_X1 U3780 ( .A1(n458), .A2(n2763), .B1(n2762), .B2(n3742), .ZN(n2192)
         );
  INV_X2 U3781 ( .A(n327), .ZN(n3744) );
  BUF_X1 U3782 ( .A(n3532), .Z(n3641) );
  BUF_X8 U3783 ( .A(n3532), .Z(n3642) );
  OR2_X2 U3784 ( .A1(n1281), .A2(n1302), .ZN(n3643) );
  OAI22_X1 U3785 ( .A1(n437), .A2(n2974), .B1(n2973), .B2(n3737), .ZN(n2410)
         );
  OAI22_X1 U3786 ( .A1(n446), .A2(n3283), .B1(n2898), .B2(n3728), .ZN(n2067)
         );
  OAI22_X1 U3787 ( .A1(n3491), .A2(n2866), .B1(n3728), .B2(n3283), .ZN(n2299)
         );
  NAND2_X1 U3788 ( .A1(n3515), .A2(n736), .ZN(n551) );
  INV_X1 U3789 ( .A(n736), .ZN(n734) );
  NAND2_X1 U3790 ( .A1(n1259), .A2(n1280), .ZN(n736) );
  XNOR2_X1 U3791 ( .A(n595), .B(n3644), .ZN(product[63]) );
  INV_X32 U3792 ( .A(n532), .ZN(n3644) );
  XNOR2_X1 U3793 ( .A(n2159), .B(n3645), .ZN(n1668) );
  XNOR2_X1 U3794 ( .A(n2607), .B(n2127), .ZN(n3645) );
  NAND2_X1 U3795 ( .A1(n1219), .A2(n1238), .ZN(n716) );
  NOR2_X1 U3796 ( .A1(n1219), .A2(n1238), .ZN(n715) );
  NAND2_X1 U3797 ( .A1(n3743), .A2(n327), .ZN(n3746) );
  INV_X1 U3798 ( .A(n3680), .ZN(n3681) );
  NAND2_X1 U3799 ( .A1(n3652), .A2(n2248), .ZN(n3646) );
  NAND2_X1 U3800 ( .A1(n3652), .A2(n2440), .ZN(n3647) );
  NAND2_X1 U3801 ( .A1(n2248), .A2(n2440), .ZN(n3648) );
  NAND3_X1 U3802 ( .A1(n3646), .A2(n3647), .A3(n3648), .ZN(n1450) );
  NAND2_X1 U3803 ( .A1(n1449), .A2(n1457), .ZN(n3649) );
  NAND2_X1 U3804 ( .A1(n1449), .A2(n1451), .ZN(n3650) );
  NAND2_X1 U3805 ( .A1(n1457), .A2(n1451), .ZN(n3651) );
  NAND3_X1 U3806 ( .A1(n3649), .A2(n3650), .A3(n3651), .ZN(n1442) );
  BUF_X1 U3807 ( .A(n2408), .Z(n3652) );
  INV_X1 U3808 ( .A(n3448), .ZN(n3680) );
  BUF_X1 U3809 ( .A(n781), .Z(n3653) );
  NAND2_X1 U3810 ( .A1(n1459), .A2(n1488), .ZN(n781) );
  OAI22_X1 U3811 ( .A1(n425), .A2(n3102), .B1(n3101), .B2(n3674), .ZN(n2542)
         );
  OAI22_X1 U3812 ( .A1(n425), .A2(n3118), .B1(n3117), .B2(n3674), .ZN(n2558)
         );
  OAI22_X1 U3813 ( .A1(n425), .A2(n3115), .B1(n3114), .B2(n3674), .ZN(n2555)
         );
  OAI22_X1 U3814 ( .A1(n425), .A2(n3111), .B1(n3110), .B2(n3674), .ZN(n2551)
         );
  OAI22_X1 U3815 ( .A1(n425), .A2(n3114), .B1(n3113), .B2(n3674), .ZN(n2554)
         );
  OAI22_X1 U3816 ( .A1(n425), .A2(n3103), .B1(n3102), .B2(n3674), .ZN(n2543)
         );
  OAI22_X1 U3817 ( .A1(n425), .A2(n3113), .B1(n3112), .B2(n3674), .ZN(n2553)
         );
  OAI22_X1 U3818 ( .A1(n425), .A2(n3097), .B1(n3674), .B2(n3290), .ZN(n2537)
         );
  OAI22_X1 U3819 ( .A1(n425), .A2(n3100), .B1(n3099), .B2(n3674), .ZN(n2540)
         );
  OAI22_X1 U3820 ( .A1(n425), .A2(n3104), .B1(n3103), .B2(n3674), .ZN(n2544)
         );
  OAI22_X1 U3821 ( .A1(n425), .A2(n3107), .B1(n3106), .B2(n3674), .ZN(n2547)
         );
  OAI22_X1 U3822 ( .A1(n437), .A2(n2972), .B1(n2971), .B2(n3737), .ZN(n2408)
         );
  INV_X1 U3823 ( .A(n3789), .ZN(n396) );
  NAND2_X1 U3824 ( .A1(n3643), .A2(n997), .ZN(n3654) );
  NAND2_X1 U3825 ( .A1(n3643), .A2(n997), .ZN(n731) );
  INV_X1 U3826 ( .A(n3539), .ZN(n3655) );
  INV_X2 U3827 ( .A(n3539), .ZN(n3657) );
  INV_X2 U3828 ( .A(n3539), .ZN(n3656) );
  NAND2_X1 U3829 ( .A1(a[6]), .A2(n3744), .ZN(n3745) );
  NAND2_X1 U3830 ( .A1(n2159), .A2(n2607), .ZN(n3658) );
  NAND2_X1 U3831 ( .A1(n2159), .A2(n2127), .ZN(n3659) );
  NAND2_X1 U3832 ( .A1(n2607), .A2(n2127), .ZN(n3660) );
  NAND3_X1 U3833 ( .A1(n3658), .A2(n3660), .A3(n3659), .ZN(n1667) );
  OR2_X1 U3834 ( .A1(n3796), .A2(n2731), .ZN(n3661) );
  OR2_X1 U3835 ( .A1(n2730), .A2(n3545), .ZN(n3662) );
  NAND2_X1 U3836 ( .A1(n3661), .A2(n3662), .ZN(n2159) );
  NOR2_X1 U3837 ( .A1(n3642), .A2(n3444), .ZN(n2127) );
  OAI22_X1 U3838 ( .A1(n419), .A2(n3165), .B1(n3164), .B2(n369), .ZN(n2607) );
  XNOR2_X1 U3839 ( .A(n469), .B(n363), .ZN(n2731) );
  XNOR2_X1 U3840 ( .A(n471), .B(n363), .ZN(n2730) );
  OAI21_X1 U3841 ( .B1(n884), .B2(n880), .A(n881), .ZN(n879) );
  OAI21_X1 U3842 ( .B1(n896), .B2(n883), .A(n884), .ZN(n882) );
  OAI22_X1 U3843 ( .A1(n3457), .A2(n2698), .B1(n2697), .B2(n3642), .ZN(n2125)
         );
  OAI22_X1 U3844 ( .A1(n3457), .A2(n2695), .B1(n2694), .B2(n3642), .ZN(n2122)
         );
  BUF_X1 U3845 ( .A(n1377), .Z(n3664) );
  NOR2_X2 U3846 ( .A1(n759), .A2(n754), .ZN(n752) );
  XOR2_X2 U3847 ( .A(n3666), .B(n1585), .Z(n1553) );
  XOR2_X2 U3848 ( .A(n3667), .B(n1553), .Z(n1551) );
  NAND2_X1 U3849 ( .A1(n1559), .A2(n1557), .ZN(n3668) );
  NAND2_X1 U3850 ( .A1(n1559), .A2(n1585), .ZN(n3669) );
  NAND2_X1 U3851 ( .A1(n1557), .A2(n1585), .ZN(n3670) );
  NAND3_X1 U3852 ( .A1(n3668), .A2(n3669), .A3(n3670), .ZN(n1552) );
  NAND2_X1 U3853 ( .A1(n1583), .A2(n1555), .ZN(n3671) );
  NAND2_X1 U3854 ( .A1(n1583), .A2(n1553), .ZN(n3672) );
  NAND2_X1 U3855 ( .A1(n1555), .A2(n1553), .ZN(n3673) );
  NAND3_X1 U3856 ( .A1(n3671), .A2(n3672), .A3(n3673), .ZN(n1550) );
  OAI22_X1 U3857 ( .A1(n3619), .A2(n3473), .B1(n3096), .B2(n3679), .ZN(n2073)
         );
  OAI22_X1 U3858 ( .A1(n3620), .A2(n3064), .B1(n3679), .B2(n3473), .ZN(n2503)
         );
  INV_X1 U3859 ( .A(n634), .ZN(n632) );
  OAI22_X1 U3860 ( .A1(n3788), .A2(n2841), .B1(n2840), .B2(n3613), .ZN(n2273)
         );
  OAI22_X1 U3861 ( .A1(n3788), .A2(n2836), .B1(n2835), .B2(n3613), .ZN(n2268)
         );
  OAI22_X1 U3862 ( .A1(n3788), .A2(n2835), .B1(n2834), .B2(n3613), .ZN(n2267)
         );
  OAI22_X1 U3863 ( .A1(n3562), .A2(n2838), .B1(n2837), .B2(n3613), .ZN(n2270)
         );
  OAI22_X1 U3864 ( .A1(n3788), .A2(n2834), .B1(n2833), .B2(n3613), .ZN(n2266)
         );
  OAI22_X1 U3865 ( .A1(n3788), .A2(n2843), .B1(n2842), .B2(n3613), .ZN(n2275)
         );
  OAI22_X1 U3866 ( .A1(n3561), .A2(n2840), .B1(n2839), .B2(n3613), .ZN(n2272)
         );
  OAI22_X1 U3867 ( .A1(n3562), .A2(n2839), .B1(n2838), .B2(n3613), .ZN(n2271)
         );
  OAI22_X1 U3868 ( .A1(n3457), .A2(n2694), .B1(n2693), .B2(n3642), .ZN(n2121)
         );
  INV_X4 U3869 ( .A(n3703), .ZN(n3674) );
  INV_X2 U3870 ( .A(n3684), .ZN(n3703) );
  INV_X1 U3871 ( .A(n3790), .ZN(n3677) );
  INV_X4 U3872 ( .A(n3676), .ZN(n3679) );
  INV_X2 U3873 ( .A(n3676), .ZN(n3678) );
  OAI22_X1 U3874 ( .A1(n431), .A2(n3039), .B1(n3038), .B2(n3656), .ZN(n2477)
         );
  OAI22_X1 U3875 ( .A1(n431), .A2(n3038), .B1(n3037), .B2(n3657), .ZN(n2476)
         );
  OAI22_X1 U3876 ( .A1(n431), .A2(n3047), .B1(n3046), .B2(n3657), .ZN(n2485)
         );
  OAI22_X1 U3877 ( .A1(n431), .A2(n3041), .B1(n3040), .B2(n3657), .ZN(n2479)
         );
  OAI22_X1 U3878 ( .A1(n431), .A2(n3034), .B1(n3033), .B2(n3656), .ZN(n2472)
         );
  OAI21_X1 U3879 ( .B1(n657), .B2(n637), .A(n638), .ZN(n636) );
  NAND2_X1 U3880 ( .A1(n690), .A2(n615), .ZN(n613) );
  AOI21_X2 U3881 ( .B1(n691), .B2(n615), .A(n616), .ZN(n614) );
  OAI22_X1 U3882 ( .A1(n3458), .A2(n2682), .B1(n2681), .B2(n3642), .ZN(n2109)
         );
  NAND2_X2 U3883 ( .A1(n1123), .A2(n1136), .ZN(n669) );
  NOR2_X1 U3884 ( .A1(n1123), .A2(n1136), .ZN(n668) );
  NOR2_X1 U3885 ( .A1(n1351), .A2(n1376), .ZN(n759) );
  OAI22_X1 U3886 ( .A1(n3457), .A2(n2693), .B1(n2692), .B2(n3642), .ZN(n2120)
         );
  AND2_X2 U3887 ( .A1(n3730), .A2(n3731), .ZN(n808) );
  OAI22_X1 U3888 ( .A1(n3457), .A2(n2699), .B1(n2698), .B2(n3642), .ZN(n2126)
         );
  OAI22_X1 U3889 ( .A1(n461), .A2(n2701), .B1(n3545), .B2(n3278), .ZN(n2129)
         );
  OAI22_X1 U3890 ( .A1(n461), .A2(n2703), .B1(n2702), .B2(n3545), .ZN(n2131)
         );
  OAI22_X1 U3891 ( .A1(n461), .A2(n2704), .B1(n2703), .B2(n3545), .ZN(n2132)
         );
  OAI22_X1 U3892 ( .A1(n461), .A2(n2708), .B1(n2707), .B2(n3545), .ZN(n2136)
         );
  OAI22_X1 U3893 ( .A1(n461), .A2(n2712), .B1(n2711), .B2(n3545), .ZN(n2140)
         );
  OAI22_X1 U3894 ( .A1(n461), .A2(n2713), .B1(n2712), .B2(n3545), .ZN(n2141)
         );
  OAI22_X1 U3895 ( .A1(n461), .A2(n2719), .B1(n2718), .B2(n3545), .ZN(n2147)
         );
  OAI22_X1 U3896 ( .A1(n461), .A2(n2717), .B1(n2716), .B2(n3545), .ZN(n2145)
         );
  OAI22_X1 U3897 ( .A1(n461), .A2(n2710), .B1(n2709), .B2(n3545), .ZN(n2138)
         );
  OAI22_X1 U3898 ( .A1(n461), .A2(n2720), .B1(n2719), .B2(n3545), .ZN(n2148)
         );
  OAI22_X1 U3899 ( .A1(n461), .A2(n2714), .B1(n2713), .B2(n3545), .ZN(n2142)
         );
  OAI22_X1 U3900 ( .A1(n3796), .A2(n2728), .B1(n2727), .B2(n3589), .ZN(n2156)
         );
  OAI22_X1 U3901 ( .A1(n461), .A2(n2716), .B1(n2715), .B2(n3545), .ZN(n2144)
         );
  OAI22_X1 U3902 ( .A1(n461), .A2(n2726), .B1(n2725), .B2(n3545), .ZN(n2154)
         );
  OAI22_X1 U3903 ( .A1(n3796), .A2(n2727), .B1(n2726), .B2(n3589), .ZN(n2155)
         );
  INV_X1 U3904 ( .A(n3411), .ZN(n684) );
  NAND2_X1 U3905 ( .A1(n686), .A2(n673), .ZN(n671) );
  BUF_X1 U3906 ( .A(n612), .Z(n3682) );
  INV_X1 U3907 ( .A(n3613), .ZN(n3683) );
  INV_X2 U3908 ( .A(n3425), .ZN(n3291) );
  BUF_X1 U3909 ( .A(n603), .Z(n3685) );
  NAND2_X1 U3910 ( .A1(n3687), .A2(a[12]), .ZN(n3688) );
  INV_X2 U3911 ( .A(n336), .ZN(n3687) );
  BUF_X1 U3912 ( .A(n775), .Z(n3691) );
  BUF_X1 U3913 ( .A(n780), .Z(n3692) );
  OAI22_X1 U3914 ( .A1(n3457), .A2(n2691), .B1(n2690), .B2(n3642), .ZN(n2118)
         );
  AOI21_X2 U3915 ( .B1(n753), .B2(n729), .A(n730), .ZN(n3780) );
  OAI22_X1 U3916 ( .A1(n446), .A2(n2890), .B1(n2889), .B2(n3729), .ZN(n2323)
         );
  NOR2_X1 U3917 ( .A1(n1551), .A2(n1581), .ZN(n3693) );
  NAND2_X1 U3918 ( .A1(n3694), .A2(n3695), .ZN(n3697) );
  NAND2_X2 U3919 ( .A1(n3696), .A2(n3697), .ZN(n3800) );
  INV_X1 U3920 ( .A(n3801), .ZN(n3694) );
  INV_X1 U3921 ( .A(n354), .ZN(n3695) );
  NOR2_X1 U3922 ( .A1(n1551), .A2(n1581), .ZN(n800) );
  OAI22_X1 U3923 ( .A1(n3712), .A2(n3127), .B1(n3126), .B2(n3674), .ZN(n2567)
         );
  INV_X4 U3924 ( .A(n3711), .ZN(n3712) );
  OAI22_X1 U3925 ( .A1(n3614), .A2(n2734), .B1(n3741), .B2(n3279), .ZN(n2163)
         );
  OAI22_X1 U3926 ( .A1(n458), .A2(n3279), .B1(n2766), .B2(n3742), .ZN(n2063)
         );
  OAI21_X1 U3927 ( .B1(n3806), .B2(n3683), .A(n3775), .ZN(n2264) );
  NAND2_X1 U3928 ( .A1(n357), .A2(n3444), .ZN(n2799) );
  OAI22_X1 U3929 ( .A1(n3704), .A2(n3280), .B1(n2799), .B2(n3581), .ZN(n2064)
         );
  NAND2_X2 U3930 ( .A1(n1351), .A2(n1376), .ZN(n760) );
  XNOR2_X2 U3931 ( .A(n3698), .B(n1491), .ZN(n1489) );
  INV_X2 U3932 ( .A(n3726), .ZN(n3728) );
  AOI21_X2 U3933 ( .B1(n878), .B2(n897), .A(n879), .ZN(n877) );
  NAND2_X1 U3934 ( .A1(a[28]), .A2(n3279), .ZN(n3701) );
  NAND2_X1 U3935 ( .A1(n3699), .A2(n3700), .ZN(n3702) );
  INV_X1 U3936 ( .A(n3279), .ZN(n3700) );
  OAI22_X1 U3937 ( .A1(n3796), .A2(n3278), .B1(n2733), .B2(n3545), .ZN(n2062)
         );
  OAI22_X1 U3938 ( .A1(n428), .A2(n3067), .B1(n3066), .B2(n3679), .ZN(n2506)
         );
  INV_X1 U3939 ( .A(n3580), .ZN(n3704) );
  INV_X4 U3940 ( .A(n3580), .ZN(n3706) );
  OAI22_X1 U3941 ( .A1(n425), .A2(n3099), .B1(n3098), .B2(n3674), .ZN(n2539)
         );
  BUF_X1 U3942 ( .A(n2345), .Z(n3707) );
  OAI22_X1 U3943 ( .A1(n446), .A2(n2896), .B1(n2895), .B2(n3729), .ZN(n2329)
         );
  NOR2_X1 U3944 ( .A1(n2022), .A2(n2029), .ZN(n934) );
  NAND2_X2 U3945 ( .A1(n2022), .A2(n2029), .ZN(n935) );
  OAI21_X1 U3946 ( .B1(n3807), .B2(n3777), .A(n363), .ZN(n2128) );
  OAI21_X1 U3947 ( .B1(n3439), .B2(n3798), .A(n3681), .ZN(n2434) );
  OAI22_X1 U3948 ( .A1(n3494), .A2(n3024), .B1(n3023), .B2(n3721), .ZN(n2461)
         );
  OAI22_X1 U3949 ( .A1(n3494), .A2(n3020), .B1(n3019), .B2(n3721), .ZN(n2457)
         );
  OAI22_X1 U3950 ( .A1(n3494), .A2(n3003), .B1(n3002), .B2(n3721), .ZN(n2440)
         );
  OAI22_X1 U3951 ( .A1(n3494), .A2(n3007), .B1(n3006), .B2(n3721), .ZN(n2444)
         );
  OAI22_X1 U3952 ( .A1(n434), .A2(n3015), .B1(n3014), .B2(n3721), .ZN(n2452)
         );
  OAI22_X1 U3953 ( .A1(n434), .A2(n3012), .B1(n3011), .B2(n3721), .ZN(n2449)
         );
  OAI22_X1 U3954 ( .A1(n434), .A2(n3013), .B1(n3012), .B2(n3721), .ZN(n2450)
         );
  OAI22_X1 U3955 ( .A1(n3494), .A2(n2998), .B1(n3721), .B2(n3287), .ZN(n2435)
         );
  OAI22_X1 U3956 ( .A1(n434), .A2(n3021), .B1(n3020), .B2(n3721), .ZN(n2458)
         );
  OAI22_X1 U3957 ( .A1(n434), .A2(n3026), .B1(n3025), .B2(n3721), .ZN(n2463)
         );
  OAI22_X1 U3958 ( .A1(n3494), .A2(n3009), .B1(n3008), .B2(n3721), .ZN(n2446)
         );
  OAI22_X1 U3959 ( .A1(n434), .A2(n3019), .B1(n3018), .B2(n3721), .ZN(n2456)
         );
  OAI22_X1 U3960 ( .A1(n434), .A2(n3022), .B1(n3021), .B2(n3721), .ZN(n2459)
         );
  OAI22_X1 U3961 ( .A1(n434), .A2(n3017), .B1(n3016), .B2(n3721), .ZN(n2454)
         );
  OAI22_X1 U3962 ( .A1(n434), .A2(n3018), .B1(n3017), .B2(n3721), .ZN(n2455)
         );
  OAI22_X1 U3963 ( .A1(n3793), .A2(n3060), .B1(n3059), .B2(n3656), .ZN(n2498)
         );
  OAI22_X1 U3964 ( .A1(n3793), .A2(n3048), .B1(n3047), .B2(n3656), .ZN(n2486)
         );
  OAI22_X1 U3965 ( .A1(n3793), .A2(n3062), .B1(n3061), .B2(n3657), .ZN(n2500)
         );
  OAI21_X1 U3966 ( .B1(n3810), .B2(n3474), .A(n333), .ZN(n2468) );
  OAI22_X1 U3967 ( .A1(n3793), .A2(n3050), .B1(n3049), .B2(n3657), .ZN(n2488)
         );
  OAI22_X1 U3968 ( .A1(n3793), .A2(n3061), .B1(n3060), .B2(n3657), .ZN(n2499)
         );
  OAI22_X1 U3969 ( .A1(n3793), .A2(n3059), .B1(n3058), .B2(n3656), .ZN(n2497)
         );
  OAI22_X1 U3970 ( .A1(n3793), .A2(n3051), .B1(n3050), .B2(n3656), .ZN(n2489)
         );
  OAI22_X1 U3971 ( .A1(n3793), .A2(n3042), .B1(n3041), .B2(n3656), .ZN(n2480)
         );
  OAI22_X1 U3972 ( .A1(n3793), .A2(n3058), .B1(n3057), .B2(n3656), .ZN(n2496)
         );
  OAI22_X1 U3973 ( .A1(n3793), .A2(n3040), .B1(n3039), .B2(n3657), .ZN(n2478)
         );
  OAI22_X1 U3974 ( .A1(n3793), .A2(n3052), .B1(n3051), .B2(n3656), .ZN(n2490)
         );
  OAI22_X1 U3975 ( .A1(n3793), .A2(n3031), .B1(n3656), .B2(n3288), .ZN(n2469)
         );
  OAI22_X1 U3976 ( .A1(n3793), .A2(n3033), .B1(n3032), .B2(n3657), .ZN(n2471)
         );
  OAI22_X1 U3977 ( .A1(n3793), .A2(n3049), .B1(n3048), .B2(n3657), .ZN(n2487)
         );
  INV_X2 U3978 ( .A(n3663), .ZN(n3710) );
  INV_X1 U3979 ( .A(n425), .ZN(n3711) );
  OAI22_X1 U3980 ( .A1(n3598), .A2(n2978), .B1(n2977), .B2(n3737), .ZN(n2414)
         );
  NOR2_X1 U3981 ( .A1(n1582), .A2(n1611), .ZN(n803) );
  OAI22_X1 U3982 ( .A1(n425), .A2(n3098), .B1(n3097), .B2(n3674), .ZN(n2538)
         );
  OAI22_X1 U3983 ( .A1(n3705), .A2(n2793), .B1(n2792), .B2(n3581), .ZN(n2223)
         );
  INV_X1 U3984 ( .A(n835), .ZN(n833) );
  OAI21_X1 U3985 ( .B1(n843), .B2(n830), .A(n831), .ZN(n829) );
  NAND2_X1 U3986 ( .A1(n1011), .A2(n3560), .ZN(n565) );
  NOR2_X2 U3987 ( .A1(n780), .A2(n3756), .ZN(n775) );
  NAND2_X1 U3988 ( .A1(n1521), .A2(n1552), .ZN(n3713) );
  NAND2_X1 U3989 ( .A1(n1521), .A2(n1523), .ZN(n3714) );
  NAND2_X1 U3990 ( .A1(n1552), .A2(n1523), .ZN(n3715) );
  NAND2_X1 U3991 ( .A1(n3716), .A2(n3717), .ZN(n3719) );
  NAND2_X2 U3992 ( .A1(n3718), .A2(n3719), .ZN(n3804) );
  INV_X1 U3993 ( .A(n3410), .ZN(n3716) );
  INV_X1 U3994 ( .A(n3708), .ZN(n3815) );
  OAI21_X1 U3995 ( .B1(n3815), .B2(n3710), .A(n3571), .ZN(n2332) );
  NAND2_X1 U3996 ( .A1(n1642), .A2(n1669), .ZN(n815) );
  XNOR2_X1 U3997 ( .A(n1405), .B(n3720), .ZN(n1403) );
  XNOR2_X1 U3998 ( .A(n1432), .B(n1407), .ZN(n3720) );
  INV_X1 U3999 ( .A(n3706), .ZN(n3816) );
  XOR2_X1 U4000 ( .A(a[10]), .B(n336), .Z(n3238) );
  NAND2_X4 U4001 ( .A1(n3242), .A2(n372), .ZN(n3722) );
  OAI22_X1 U4002 ( .A1(n434), .A2(n3006), .B1(n3721), .B2(n3005), .ZN(n2443)
         );
  INV_X1 U4003 ( .A(n3548), .ZN(n855) );
  INV_X1 U4004 ( .A(n887), .ZN(n885) );
  INV_X1 U4005 ( .A(n3692), .ZN(n1005) );
  OAI21_X1 U4006 ( .B1(n3814), .B2(n3809), .A(n3425), .ZN(n2570) );
  NAND2_X1 U4007 ( .A1(n809), .A2(n817), .ZN(n807) );
  OAI21_X1 U4008 ( .B1(n3816), .B2(n3800), .A(n357), .ZN(n2196) );
  OAI22_X1 U4009 ( .A1(n3457), .A2(n2696), .B1(n2695), .B2(n3642), .ZN(n2123)
         );
  INV_X1 U4010 ( .A(n3726), .ZN(n3727) );
  INV_X4 U4011 ( .A(n3726), .ZN(n3729) );
  OAI22_X1 U4012 ( .A1(n434), .A2(n3005), .B1(n3004), .B2(n3721), .ZN(n2442)
         );
  NAND2_X1 U4013 ( .A1(n809), .A2(n818), .ZN(n3730) );
  INV_X1 U4014 ( .A(n810), .ZN(n3731) );
  OAI21_X1 U4015 ( .B1(n782), .B2(n3692), .A(n3653), .ZN(n779) );
  NOR2_X2 U4016 ( .A1(n784), .A2(n765), .ZN(n763) );
  INV_X2 U4017 ( .A(n387), .ZN(n3734) );
  INV_X8 U4018 ( .A(n3811), .ZN(n425) );
  NAND2_X1 U4019 ( .A1(n1491), .A2(n3440), .ZN(n3738) );
  NAND2_X1 U4020 ( .A1(n1491), .A2(n1493), .ZN(n3739) );
  NAND2_X1 U4021 ( .A1(n3440), .A2(n1493), .ZN(n3740) );
  NAND3_X1 U4022 ( .A1(n3738), .A2(n3740), .A3(n3739), .ZN(n1488) );
  NOR2_X2 U4023 ( .A1(n1459), .A2(n1488), .ZN(n780) );
  INV_X1 U4024 ( .A(n3792), .ZN(n408) );
  OAI21_X1 U4025 ( .B1(n3690), .B2(n3791), .A(n366), .ZN(n3817) );
  OAI21_X1 U4026 ( .B1(n3803), .B2(n3789), .A(n348), .ZN(n2298) );
  OAI21_X1 U4027 ( .B1(n3725), .B2(n3804), .A(n3603), .ZN(n2366) );
  OAI22_X1 U4028 ( .A1(n3457), .A2(n3575), .B1(n2700), .B2(n3642), .ZN(n2061)
         );
  OAI21_X1 U4029 ( .B1(n3811), .B2(n3703), .A(n327), .ZN(n2536) );
  OAI21_X1 U4030 ( .B1(n816), .B2(n814), .A(n3560), .ZN(n813) );
  INV_X1 U4031 ( .A(n814), .ZN(n1011) );
  OAI21_X1 U4032 ( .B1(n3805), .B2(n3733), .A(n339), .ZN(n2400) );
  NAND2_X1 U4033 ( .A1(n885), .A2(n888), .ZN(n577) );
  INV_X1 U4034 ( .A(n877), .ZN(n876) );
  NAND2_X1 U4035 ( .A1(n885), .A2(n892), .ZN(n883) );
  OAI21_X1 U4036 ( .B1(n3802), .B2(n3790), .A(n3795), .ZN(n2502) );
  OAI22_X1 U4037 ( .A1(n440), .A2(n2949), .B1(n2948), .B2(n3626), .ZN(n2384)
         );
  OAI21_X1 U4038 ( .B1(n3808), .B2(n3792), .A(n360), .ZN(n2162) );
  XNOR2_X2 U4039 ( .A(n3282), .B(a[22]), .ZN(n3747) );
  BUF_X1 U4040 ( .A(n3577), .Z(n3748) );
  BUF_X1 U4041 ( .A(n829), .Z(n3749) );
  OAI21_X1 U4042 ( .B1(n728), .B2(n688), .A(n689), .ZN(n687) );
  XOR2_X1 U4043 ( .A(n2509), .B(n2285), .Z(n3750) );
  XOR2_X1 U4044 ( .A(n3755), .B(n3750), .Z(n1604) );
  NAND2_X1 U4045 ( .A1(n3755), .A2(n2509), .ZN(n3751) );
  NAND2_X1 U4046 ( .A1(n3755), .A2(n2285), .ZN(n3752) );
  NAND2_X1 U4047 ( .A1(n2509), .A2(n2285), .ZN(n3753) );
  NAND3_X1 U4048 ( .A1(n3751), .A2(n3753), .A3(n3752), .ZN(n1603) );
  BUF_X2 U4049 ( .A(n2253), .Z(n3755) );
  OAI22_X1 U4050 ( .A1(n3619), .A2(n3070), .B1(n3069), .B2(n3678), .ZN(n2509)
         );
  NAND2_X1 U4051 ( .A1(n1018), .A2(n862), .ZN(n572) );
  NAND2_X1 U4052 ( .A1(n859), .A2(n867), .ZN(n857) );
  XNOR2_X1 U4053 ( .A(n863), .B(n572), .ZN(product[23]) );
  NAND2_X1 U4054 ( .A1(n1002), .A2(n770), .ZN(n556) );
  NAND2_X1 U4055 ( .A1(n1377), .A2(n1402), .ZN(n770) );
  XNOR2_X1 U4056 ( .A(n771), .B(n556), .ZN(product[39]) );
  XOR2_X1 U4057 ( .A(n774), .B(n557), .Z(product[38]) );
  OAI21_X1 U4058 ( .B1(n855), .B2(n842), .A(n3442), .ZN(n841) );
  NAND2_X1 U4059 ( .A1(n1004), .A2(n778), .ZN(n558) );
  NAND2_X1 U4060 ( .A1(n3785), .A2(n789), .ZN(n560) );
  NAND2_X1 U4061 ( .A1(n791), .A2(n794), .ZN(n561) );
  INV_X1 U4062 ( .A(n794), .ZN(n792) );
  XOR2_X1 U4063 ( .A(n1447), .B(n1472), .Z(n3757) );
  XOR2_X1 U4064 ( .A(n3757), .B(n1470), .Z(n1439) );
  XOR2_X1 U4065 ( .A(n1466), .B(n1441), .Z(n3758) );
  XOR2_X1 U4066 ( .A(n3758), .B(n1439), .Z(n1435) );
  NAND2_X1 U4067 ( .A1(n1447), .A2(n1472), .ZN(n3759) );
  NAND2_X1 U4068 ( .A1(n1447), .A2(n1470), .ZN(n3760) );
  NAND2_X1 U4069 ( .A1(n1472), .A2(n1470), .ZN(n3761) );
  NAND3_X1 U4070 ( .A1(n3759), .A2(n3760), .A3(n3761), .ZN(n1438) );
  NAND2_X1 U4071 ( .A1(n1466), .A2(n1441), .ZN(n3762) );
  NAND2_X1 U4072 ( .A1(n1466), .A2(n1439), .ZN(n3763) );
  NAND2_X1 U4073 ( .A1(n1441), .A2(n1439), .ZN(n3764) );
  NAND3_X1 U4074 ( .A1(n3762), .A2(n3763), .A3(n3764), .ZN(n1434) );
  XOR2_X1 U4075 ( .A(n2313), .B(n2345), .Z(n3765) );
  XOR2_X1 U4076 ( .A(n2249), .B(n3765), .Z(n1477) );
  NAND2_X1 U4077 ( .A1(n2249), .A2(n2313), .ZN(n3766) );
  NAND2_X1 U4078 ( .A1(n2249), .A2(n3707), .ZN(n3767) );
  NAND2_X1 U4079 ( .A1(n2313), .A2(n3707), .ZN(n3768) );
  NAND3_X1 U4080 ( .A1(n3766), .A2(n3768), .A3(n3767), .ZN(n1476) );
  BUF_X1 U4081 ( .A(n749), .Z(n3769) );
  OAI22_X1 U4082 ( .A1(n446), .A2(n2880), .B1(n2879), .B2(n3729), .ZN(n2313)
         );
  OAI22_X1 U4083 ( .A1(n443), .A2(n2911), .B1(n2910), .B2(n393), .ZN(n2345) );
  AOI21_X1 U4084 ( .B1(n749), .B2(n999), .A(n746), .ZN(n744) );
  NAND2_X1 U4085 ( .A1(n786), .A2(n798), .ZN(n784) );
  NAND2_X1 U4086 ( .A1(n1405), .A2(n1432), .ZN(n3770) );
  NAND2_X1 U4087 ( .A1(n1405), .A2(n1407), .ZN(n3771) );
  NAND2_X1 U4088 ( .A1(n1432), .A2(n1407), .ZN(n3772) );
  NAND3_X1 U4089 ( .A1(n3770), .A2(n3772), .A3(n3771), .ZN(n1402) );
  INV_X1 U4090 ( .A(n3799), .ZN(n3779) );
  INV_X1 U4091 ( .A(n754), .ZN(n1000) );
  NAND2_X1 U4092 ( .A1(n1327), .A2(n1350), .ZN(n755) );
  NOR2_X2 U4093 ( .A1(n1327), .A2(n1350), .ZN(n754) );
  OR2_X1 U4094 ( .A1(n1551), .A2(n1581), .ZN(n3773) );
  AOI21_X1 U4095 ( .B1(n826), .B2(n817), .A(n3564), .ZN(n816) );
  INV_X1 U4096 ( .A(n819), .ZN(n1012) );
  NOR2_X2 U4097 ( .A1(n1670), .A2(n1697), .ZN(n819) );
  NOR2_X1 U4098 ( .A1(n803), .A2(n3693), .ZN(n798) );
  OAI21_X1 U4099 ( .B1(n3780), .B2(n613), .A(n614), .ZN(n612) );
  BUF_X1 U4100 ( .A(n776), .Z(n3774) );
  OAI21_X1 U4101 ( .B1(n777), .B2(n781), .A(n778), .ZN(n776) );
  INV_X1 U4102 ( .A(n3446), .ZN(n1018) );
  OAI21_X1 U4103 ( .B1(n3475), .B2(n865), .A(n862), .ZN(n860) );
  NAND2_X1 U4104 ( .A1(n1820), .A2(n1841), .ZN(n862) );
  OAI22_X1 U4105 ( .A1(n3561), .A2(n2833), .B1(n3613), .B2(n3282), .ZN(n2265)
         );
  INV_X16 U4106 ( .A(a[0]), .ZN(n369) );
  INV_X1 U4107 ( .A(n687), .ZN(n685) );
  AOI21_X2 U4108 ( .B1(n687), .B2(n673), .A(n676), .ZN(n672) );
  OAI22_X1 U4109 ( .A1(n3441), .A2(n2816), .B1(n2815), .B2(n402), .ZN(n2247)
         );
  OAI22_X1 U4110 ( .A1(n3778), .A2(n2813), .B1(n2812), .B2(n402), .ZN(n2244)
         );
  OAI22_X1 U4111 ( .A1(n3441), .A2(n2804), .B1(n2803), .B2(n402), .ZN(n2235)
         );
  OAI22_X1 U4112 ( .A1(n3778), .A2(n2814), .B1(n2813), .B2(n402), .ZN(n2245)
         );
  OAI22_X1 U4113 ( .A1(n3778), .A2(n2809), .B1(n2808), .B2(n402), .ZN(n2240)
         );
  OAI22_X1 U4114 ( .A1(n3778), .A2(n2810), .B1(n2809), .B2(n402), .ZN(n2241)
         );
  OAI22_X1 U4115 ( .A1(n3778), .A2(n2812), .B1(n2811), .B2(n402), .ZN(n2243)
         );
  OAI22_X1 U4116 ( .A1(n3778), .A2(n2806), .B1(n2805), .B2(n402), .ZN(n2237)
         );
  OAI22_X1 U4117 ( .A1(n3508), .A2(n2815), .B1(n2814), .B2(n402), .ZN(n2246)
         );
  OAI22_X1 U4118 ( .A1(n3779), .A2(n3281), .B1(n2832), .B2(n402), .ZN(n2065)
         );
  OAI22_X1 U4119 ( .A1(n3779), .A2(n2817), .B1(n2816), .B2(n402), .ZN(n2248)
         );
  OAI22_X1 U4120 ( .A1(n3778), .A2(n2805), .B1(n2804), .B2(n402), .ZN(n2236)
         );
  INV_X2 U4121 ( .A(n3282), .ZN(n3775) );
  AOI21_X1 U4122 ( .B1(n783), .B2(n3691), .A(n3774), .ZN(n774) );
  OAI22_X1 U4123 ( .A1(n3441), .A2(n2808), .B1(n2807), .B2(n402), .ZN(n2239)
         );
  OAI22_X1 U4124 ( .A1(n3441), .A2(n2803), .B1(n2802), .B2(n402), .ZN(n2234)
         );
  OAI22_X1 U4125 ( .A1(n3778), .A2(n2800), .B1(n402), .B2(n3281), .ZN(n2231)
         );
  OAI22_X1 U4126 ( .A1(n3778), .A2(n2801), .B1(n2800), .B2(n402), .ZN(n2232)
         );
  OAI22_X1 U4127 ( .A1(n3778), .A2(n2807), .B1(n2806), .B2(n402), .ZN(n2238)
         );
  OAI22_X1 U4128 ( .A1(n3778), .A2(n2802), .B1(n2801), .B2(n402), .ZN(n2233)
         );
  OAI22_X1 U4129 ( .A1(n2811), .A2(n3779), .B1(n2810), .B2(n402), .ZN(n2242)
         );
  OAI22_X1 U4130 ( .A1(n3778), .A2(n2831), .B1(n2830), .B2(n402), .ZN(n2262)
         );
  NOR2_X2 U4131 ( .A1(n1642), .A2(n1669), .ZN(n814) );
  NOR2_X1 U4132 ( .A1(n1918), .A2(n1933), .ZN(n887) );
  NAND2_X2 U4133 ( .A1(n1918), .A2(n1933), .ZN(n888) );
  NAND2_X1 U4134 ( .A1(n1489), .A2(n3409), .ZN(n789) );
  OAI21_X1 U4135 ( .B1(n3605), .B2(n815), .A(n812), .ZN(n810) );
  NAND2_X1 U4136 ( .A1(n1612), .A2(n1641), .ZN(n812) );
  INV_X4 U4137 ( .A(n360), .ZN(n3279) );
  AND2_X2 U4138 ( .A1(n3786), .A2(n3787), .ZN(n785) );
  OAI22_X1 U4139 ( .A1(n3509), .A2(n2818), .B1(n2817), .B2(n402), .ZN(n2249)
         );
  OAI22_X1 U4140 ( .A1(n3509), .A2(n2820), .B1(n2819), .B2(n402), .ZN(n2251)
         );
  OAI22_X1 U4141 ( .A1(n3509), .A2(n2822), .B1(n2821), .B2(n402), .ZN(n2253)
         );
  OAI22_X1 U4142 ( .A1(n3471), .A2(n2827), .B1(n2826), .B2(n402), .ZN(n2258)
         );
  OAI22_X1 U4143 ( .A1(n2830), .A2(n3508), .B1(n2829), .B2(n402), .ZN(n2261)
         );
  OAI22_X1 U4144 ( .A1(n3509), .A2(n2823), .B1(n2822), .B2(n402), .ZN(n2254)
         );
  OAI22_X1 U4145 ( .A1(n3509), .A2(n2826), .B1(n2825), .B2(n402), .ZN(n2257)
         );
  OAI22_X1 U4146 ( .A1(n2819), .A2(n3508), .B1(n2818), .B2(n402), .ZN(n2250)
         );
  INV_X4 U4147 ( .A(n351), .ZN(n3282) );
  AOI21_X1 U4148 ( .B1(n753), .B2(n729), .A(n730), .ZN(n728) );
  OAI21_X1 U4149 ( .B1(n731), .B2(n748), .A(n732), .ZN(n730) );
  AOI21_X2 U4150 ( .B1(n997), .B2(n3665), .A(n734), .ZN(n732) );
  NAND2_X1 U4151 ( .A1(n844), .A2(n847), .ZN(n570) );
  NAND2_X2 U4152 ( .A1(n844), .A2(n851), .ZN(n842) );
  NOR2_X2 U4153 ( .A1(n1774), .A2(n1797), .ZN(n846) );
  NAND2_X1 U4154 ( .A1(n1774), .A2(n1797), .ZN(n847) );
  NAND2_X2 U4155 ( .A1(n1670), .A2(n1697), .ZN(n820) );
  NOR2_X1 U4156 ( .A1(n3664), .A2(n1402), .ZN(n3782) );
  NAND2_X2 U4157 ( .A1(n3604), .A2(n3576), .ZN(n830) );
  AOI21_X1 U4158 ( .B1(n841), .B2(n3576), .A(n838), .ZN(n836) );
  NAND2_X1 U4159 ( .A1(n3576), .A2(n840), .ZN(n569) );
  OAI22_X1 U4160 ( .A1(n3509), .A2(n2828), .B1(n2827), .B2(n402), .ZN(n2259)
         );
  NAND2_X2 U4161 ( .A1(n1724), .A2(n1749), .ZN(n835) );
  NAND2_X1 U4162 ( .A1(n1009), .A2(n3748), .ZN(n563) );
  OAI21_X1 U4163 ( .B1(n805), .B2(n803), .A(n3748), .ZN(n802) );
  NAND2_X1 U4164 ( .A1(n1582), .A2(n1611), .ZN(n804) );
  BUF_X1 U4165 ( .A(n3635), .Z(n3783) );
  OAI22_X1 U4166 ( .A1(n3565), .A2(n2824), .B1(n2823), .B2(n402), .ZN(n2255)
         );
  AOI21_X1 U4167 ( .B1(n3548), .B2(n828), .A(n3749), .ZN(n3784) );
  OAI21_X2 U4168 ( .B1(n827), .B2(n807), .A(n808), .ZN(n806) );
  AOI21_X2 U4169 ( .B1(n856), .B2(n828), .A(n829), .ZN(n827) );
  INV_X1 U4170 ( .A(n3754), .ZN(n791) );
  NAND2_X1 U4171 ( .A1(n1431), .A2(n1458), .ZN(n778) );
  INV_X1 U4172 ( .A(n3537), .ZN(n1004) );
  OAI21_X1 U4173 ( .B1(n3799), .B2(n3747), .A(n354), .ZN(n2230) );
  NAND2_X1 U4174 ( .A1(n1005), .A2(n3653), .ZN(n559) );
  INV_X1 U4175 ( .A(n3497), .ZN(n1003) );
  OAI21_X1 U4176 ( .B1(n774), .B2(n3497), .A(n773), .ZN(n771) );
  NOR2_X2 U4177 ( .A1(n769), .A2(n772), .ZN(n767) );
  NOR2_X2 U4178 ( .A1(n1403), .A2(n1430), .ZN(n772) );
  NAND2_X2 U4179 ( .A1(n1403), .A2(n1430), .ZN(n773) );
  INV_X1 U4180 ( .A(n3780), .ZN(n726) );
  OAI22_X1 U4181 ( .A1(n3788), .A2(n2859), .B1(n2858), .B2(n3613), .ZN(n2291)
         );
  OAI22_X1 U4182 ( .A1(n3561), .A2(n2844), .B1(n2843), .B2(n3613), .ZN(n2276)
         );
  OAI22_X1 U4183 ( .A1(n3562), .A2(n2842), .B1(n2841), .B2(n3613), .ZN(n2274)
         );
  OAI22_X1 U4184 ( .A1(n3561), .A2(n2837), .B1(n2836), .B2(n3613), .ZN(n2269)
         );
  OAI22_X1 U4185 ( .A1(n3562), .A2(n2858), .B1(n2857), .B2(n3613), .ZN(n2290)
         );
  OAI22_X1 U4186 ( .A1(n3561), .A2(n2862), .B1(n2861), .B2(n3613), .ZN(n2294)
         );
  OAI22_X1 U4187 ( .A1(n3562), .A2(n2848), .B1(n2847), .B2(n3613), .ZN(n2280)
         );
  OAI22_X1 U4188 ( .A1(n3561), .A2(n2847), .B1(n2846), .B2(n3613), .ZN(n2279)
         );
  OAI22_X1 U4189 ( .A1(n449), .A2(n2853), .B1(n2852), .B2(n3613), .ZN(n2285)
         );
  OAI22_X1 U4190 ( .A1(n3562), .A2(n2857), .B1(n2856), .B2(n3613), .ZN(n2289)
         );
  OAI22_X1 U4191 ( .A1(n3562), .A2(n2851), .B1(n2850), .B2(n3613), .ZN(n2283)
         );
  OAI22_X1 U4192 ( .A1(n3562), .A2(n2864), .B1(n2863), .B2(n3613), .ZN(n2296)
         );
  OAI22_X1 U4193 ( .A1(n3561), .A2(n2845), .B1(n2844), .B2(n3613), .ZN(n2277)
         );
  OAI22_X1 U4194 ( .A1(n3561), .A2(n3282), .B1(n2865), .B2(n3613), .ZN(n2066)
         );
  OAI22_X1 U4195 ( .A1(n3788), .A2(n2855), .B1(n2854), .B2(n3613), .ZN(n2287)
         );
  OAI22_X1 U4196 ( .A1(n449), .A2(n2860), .B1(n2859), .B2(n3613), .ZN(n2292)
         );
  OAI22_X1 U4197 ( .A1(n3562), .A2(n2861), .B1(n2860), .B2(n3613), .ZN(n2293)
         );
  OAI22_X1 U4198 ( .A1(n3561), .A2(n2850), .B1(n2849), .B2(n3613), .ZN(n2282)
         );
  OAI22_X1 U4199 ( .A1(n3562), .A2(n2863), .B1(n2862), .B2(n3613), .ZN(n2295)
         );
  OAI22_X1 U4200 ( .A1(n3561), .A2(n2849), .B1(n2848), .B2(n3613), .ZN(n2281)
         );
  OAI22_X1 U4201 ( .A1(n3562), .A2(n2846), .B1(n2845), .B2(n3613), .ZN(n2278)
         );
  OAI22_X1 U4202 ( .A1(n3561), .A2(n2856), .B1(n2855), .B2(n3613), .ZN(n2288)
         );
  OAI22_X1 U4203 ( .A1(n449), .A2(n2852), .B1(n2851), .B2(n3612), .ZN(n2284)
         );
  OAI22_X1 U4204 ( .A1(n3794), .A2(n3056), .B1(n3055), .B2(n3657), .ZN(n2494)
         );
  OAI22_X1 U4205 ( .A1(n3794), .A2(n3288), .B1(n3063), .B2(n3656), .ZN(n2072)
         );
  OAI22_X1 U4206 ( .A1(n3794), .A2(n3036), .B1(n3035), .B2(n3656), .ZN(n2474)
         );
  OAI22_X1 U4207 ( .A1(n3794), .A2(n3054), .B1(n3053), .B2(n3657), .ZN(n2492)
         );
  OAI22_X1 U4208 ( .A1(n3794), .A2(n3055), .B1(n3054), .B2(n3657), .ZN(n2493)
         );
  OAI22_X1 U4209 ( .A1(n3794), .A2(n3057), .B1(n3056), .B2(n3656), .ZN(n2495)
         );
  OAI22_X1 U4210 ( .A1(n3794), .A2(n3045), .B1(n3044), .B2(n3657), .ZN(n2483)
         );
  OAI22_X1 U4211 ( .A1(n3794), .A2(n3044), .B1(n3043), .B2(n3656), .ZN(n2482)
         );
  OAI22_X1 U4212 ( .A1(n3794), .A2(n3046), .B1(n3045), .B2(n3656), .ZN(n2484)
         );
  OAI22_X1 U4213 ( .A1(n3794), .A2(n3032), .B1(n3031), .B2(n3656), .ZN(n2470)
         );
  OAI22_X1 U4214 ( .A1(n3794), .A2(n3053), .B1(n3052), .B2(n3657), .ZN(n2491)
         );
  OAI22_X1 U4215 ( .A1(n3794), .A2(n3035), .B1(n3034), .B2(n3657), .ZN(n2473)
         );
  OAI22_X1 U4216 ( .A1(n3794), .A2(n3037), .B1(n3036), .B2(n3657), .ZN(n2475)
         );
  OAI22_X1 U4217 ( .A1(n3794), .A2(n3043), .B1(n3042), .B2(n3656), .ZN(n2481)
         );
  INV_X1 U4218 ( .A(n3784), .ZN(n826) );
  XOR2_X1 U4219 ( .A(n682), .B(n545), .Z(product[50]) );
  OAI21_X2 U4220 ( .B1(n682), .B2(n680), .A(n681), .ZN(n679) );
  OR2_X1 U4221 ( .A1(n1489), .A2(n3409), .ZN(n3785) );
  NAND2_X1 U4222 ( .A1(n799), .A2(n786), .ZN(n3786) );
  INV_X1 U4223 ( .A(n787), .ZN(n3787) );
  AOI21_X2 U4224 ( .B1(n776), .B2(n767), .A(n768), .ZN(n766) );
  OAI21_X1 U4225 ( .B1(n3781), .B2(n773), .A(n770), .ZN(n768) );
  OAI22_X1 U4226 ( .A1(n437), .A2(n2983), .B1(n2982), .B2(n3736), .ZN(n2419)
         );
  INV_X1 U4227 ( .A(n3783), .ZN(n797) );
  OAI22_X1 U4228 ( .A1(n461), .A2(n2702), .B1(n2701), .B2(n3545), .ZN(n2130)
         );
  OAI22_X1 U4229 ( .A1(n461), .A2(n2705), .B1(n2704), .B2(n3545), .ZN(n2133)
         );
  OAI22_X1 U4230 ( .A1(n461), .A2(n2709), .B1(n2708), .B2(n3545), .ZN(n2137)
         );
  OAI22_X1 U4231 ( .A1(n461), .A2(n2706), .B1(n2705), .B2(n3545), .ZN(n2134)
         );
  OAI22_X1 U4232 ( .A1(n461), .A2(n2707), .B1(n2706), .B2(n3545), .ZN(n2135)
         );
  OAI22_X1 U4233 ( .A1(n461), .A2(n2711), .B1(n2710), .B2(n3545), .ZN(n2139)
         );
  OAI22_X1 U4234 ( .A1(n461), .A2(n2715), .B1(n2714), .B2(n3545), .ZN(n2143)
         );
  OAI22_X1 U4235 ( .A1(n461), .A2(n2721), .B1(n2720), .B2(n3545), .ZN(n2149)
         );
  OAI22_X1 U4236 ( .A1(n461), .A2(n2718), .B1(n2717), .B2(n3545), .ZN(n2146)
         );
  OAI22_X1 U4237 ( .A1(n461), .A2(n2724), .B1(n2723), .B2(n3545), .ZN(n2152)
         );
  OAI22_X1 U4238 ( .A1(n3796), .A2(n2725), .B1(n2724), .B2(n3589), .ZN(n2153)
         );
  OAI22_X1 U4239 ( .A1(n461), .A2(n2723), .B1(n2722), .B2(n3545), .ZN(n2151)
         );
  OAI22_X1 U4240 ( .A1(n461), .A2(n2730), .B1(n2729), .B2(n3545), .ZN(n2158)
         );
  OAI22_X1 U4241 ( .A1(n461), .A2(n2732), .B1(n2731), .B2(n3545), .ZN(n2160)
         );
  OAI22_X1 U4242 ( .A1(n3796), .A2(n2722), .B1(n2721), .B2(n3589), .ZN(n2150)
         );
  OAI22_X1 U4243 ( .A1(n461), .A2(n2729), .B1(n2728), .B2(n3589), .ZN(n2157)
         );
  XNOR2_X1 U4244 ( .A(n662), .B(n541), .ZN(product[54]) );
  INV_X1 U4245 ( .A(n683), .ZN(n682) );
  XNOR2_X1 U4246 ( .A(n737), .B(n551), .ZN(product[44]) );
  INV_X1 U4247 ( .A(n3289), .ZN(n3795) );
  XNOR2_X1 U4248 ( .A(n650), .B(n539), .ZN(product[56]) );
  AOI21_X1 U4249 ( .B1(n603), .B2(n980), .A(n600), .ZN(n3797) );
  OAI22_X1 U4250 ( .A1(n3788), .A2(n2854), .B1(n2853), .B2(n3613), .ZN(n2286)
         );
  OAI21_X1 U4251 ( .B1(n788), .B2(n794), .A(n789), .ZN(n787) );
  NOR2_X2 U4252 ( .A1(n1489), .A2(n1518), .ZN(n788) );
  OAI21_X2 U4253 ( .B1(n531), .B2(n671), .A(n672), .ZN(n670) );
  OAI22_X1 U4254 ( .A1(n446), .A2(n2883), .B1(n2882), .B2(n3728), .ZN(n2316)
         );
  OAI22_X1 U4255 ( .A1(n3598), .A2(n2976), .B1(n2975), .B2(n3736), .ZN(n2412)
         );
  INV_X4 U4256 ( .A(n3807), .ZN(n461) );
  OAI22_X1 U4257 ( .A1(n3457), .A2(n2697), .B1(n2696), .B2(n3642), .ZN(n2124)
         );
  OAI21_X2 U4258 ( .B1(n630), .B2(n624), .A(n625), .ZN(n623) );
  XOR2_X1 U4259 ( .A(n630), .B(n537), .Z(product[58]) );
  AOI21_X2 U4260 ( .B1(n683), .B2(n631), .A(n632), .ZN(n630) );
  OAI21_X2 U4261 ( .B1(n701), .B2(n699), .A(n700), .ZN(n698) );
  XOR2_X1 U4262 ( .A(n701), .B(n547), .Z(product[48]) );
  AOI21_X2 U4263 ( .B1(n706), .B2(n994), .A(n703), .ZN(n701) );
  AOI21_X2 U4264 ( .B1(n670), .B2(n989), .A(n667), .ZN(n665) );
  INV_X8 U4265 ( .A(n3710), .ZN(n393) );
  XNOR2_X1 U4266 ( .A(n3769), .B(n553), .ZN(product[42]) );
  OAI21_X1 U4267 ( .B1(n744), .B2(n738), .A(n739), .ZN(n737) );
  XOR2_X1 U4268 ( .A(n744), .B(n552), .Z(product[43]) );
  XNOR2_X1 U4269 ( .A(n643), .B(n538), .ZN(product[57]) );
  OAI21_X2 U4270 ( .B1(n785), .B2(n765), .A(n766), .ZN(n764) );
  XNOR2_X1 U4271 ( .A(n3582), .B(n548), .ZN(product[47]) );
  XNOR2_X1 U4272 ( .A(n761), .B(n555), .ZN(product[40]) );
  OAI21_X1 U4273 ( .B1(n724), .B2(n718), .A(n719), .ZN(n717) );
  XOR2_X1 U4274 ( .A(n724), .B(n550), .Z(product[45]) );
  AOI21_X1 U4275 ( .B1(n761), .B2(n757), .A(n758), .ZN(n756) );
  AOI21_X1 U4276 ( .B1(n761), .B2(n611), .A(n3682), .ZN(n610) );
  AOI21_X2 U4277 ( .B1(n761), .B2(n725), .A(n726), .ZN(n724) );
  INV_X1 U4278 ( .A(n422), .ZN(n3814) );
  OAI22_X1 U4279 ( .A1(n422), .A2(n3131), .B1(n3130), .B2(n372), .ZN(n2572) );
  XNOR2_X1 U4280 ( .A(n3685), .B(n534), .ZN(product[61]) );
  XOR2_X1 U4281 ( .A(n665), .B(n542), .Z(product[53]) );
  OAI21_X1 U4282 ( .B1(n665), .B2(n663), .A(n664), .ZN(n662) );
  AOI21_X2 U4283 ( .B1(n670), .B2(n654), .A(n655), .ZN(n653) );
  AND2_X2 U4284 ( .A1(n3241), .A2(n375), .ZN(n3811) );
  XNOR2_X1 U4285 ( .A(n670), .B(n543), .ZN(product[52]) );
  OAI21_X1 U4286 ( .B1(n653), .B2(n644), .A(n645), .ZN(n643) );
  OAI21_X1 U4287 ( .B1(n653), .B2(n651), .A(n652), .ZN(n650) );
  XOR2_X1 U4288 ( .A(n653), .B(n540), .Z(product[55]) );
  INV_X1 U4289 ( .A(n531), .ZN(n761) );
  OAI21_X1 U4290 ( .B1(n750), .B2(n531), .A(n751), .ZN(n749) );
  OAI21_X1 U4291 ( .B1(n531), .B2(n684), .A(n685), .ZN(n683) );
  OAI21_X1 U4292 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  XOR2_X1 U4293 ( .A(n3797), .B(n533), .Z(product[62]) );
  INV_X2 U4294 ( .A(n594), .ZN(product[1]) );
  INV_X2 U4295 ( .A(n699), .ZN(n993) );
  INV_X2 U4296 ( .A(n680), .ZN(n991) );
  INV_X2 U4297 ( .A(n677), .ZN(n990) );
  INV_X2 U4298 ( .A(n663), .ZN(n988) );
  INV_X2 U4299 ( .A(n660), .ZN(n987) );
  INV_X2 U4300 ( .A(n651), .ZN(n986) );
  INV_X2 U4301 ( .A(n648), .ZN(n985) );
  INV_X2 U4302 ( .A(n596), .ZN(n979) );
  INV_X2 U4303 ( .A(n978), .ZN(n976) );
  INV_X2 U4304 ( .A(n975), .ZN(n973) );
  INV_X2 U4305 ( .A(n967), .ZN(n965) );
  INV_X2 U4306 ( .A(n959), .ZN(n957) );
  INV_X2 U4307 ( .A(n955), .ZN(n954) );
  INV_X2 U4308 ( .A(n953), .ZN(n951) );
  INV_X2 U4309 ( .A(n948), .ZN(n946) );
  INV_X2 U4310 ( .A(n941), .ZN(n939) );
  INV_X2 U4311 ( .A(n937), .ZN(n936) );
  INV_X2 U4312 ( .A(n935), .ZN(n933) );
  INV_X2 U4313 ( .A(n930), .ZN(n928) );
  INV_X2 U4314 ( .A(n924), .ZN(n923) );
  INV_X2 U4315 ( .A(n915), .ZN(n914) );
  INV_X2 U4316 ( .A(n913), .ZN(n911) );
  INV_X2 U4317 ( .A(n903), .ZN(n901) );
  INV_X2 U4318 ( .A(n897), .ZN(n896) );
  INV_X2 U4319 ( .A(n891), .ZN(n893) );
  INV_X2 U4320 ( .A(n888), .ZN(n886) );
  INV_X2 U4321 ( .A(n875), .ZN(n873) );
  INV_X2 U4322 ( .A(n783), .ZN(n782) );
  INV_X2 U4323 ( .A(n760), .ZN(n758) );
  INV_X2 U4324 ( .A(n752), .ZN(n750) );
  INV_X2 U4325 ( .A(n748), .ZN(n746) );
  INV_X2 U4326 ( .A(n747), .ZN(n999) );
  INV_X2 U4327 ( .A(n719), .ZN(n721) );
  INV_X2 U4328 ( .A(n715), .ZN(n995) );
  INV_X2 U4329 ( .A(n705), .ZN(n703) );
  INV_X2 U4330 ( .A(n704), .ZN(n994) );
  INV_X2 U4331 ( .A(n691), .ZN(n689) );
  INV_X2 U4332 ( .A(n669), .ZN(n667) );
  INV_X2 U4333 ( .A(n668), .ZN(n989) );
  INV_X2 U4334 ( .A(n657), .ZN(n655) );
  INV_X2 U4335 ( .A(n656), .ZN(n654) );
  INV_X2 U4336 ( .A(n647), .ZN(n645) );
  INV_X2 U4337 ( .A(n646), .ZN(n644) );
  INV_X2 U4338 ( .A(n642), .ZN(n640) );
  INV_X2 U4339 ( .A(n641), .ZN(n984) );
  INV_X2 U4340 ( .A(n633), .ZN(n631) );
  INV_X2 U4341 ( .A(n625), .ZN(n627) );
  INV_X2 U4342 ( .A(n624), .ZN(n983) );
  INV_X2 U4343 ( .A(n622), .ZN(n620) );
  INV_X2 U4344 ( .A(n621), .ZN(n982) );
  INV_X2 U4345 ( .A(n609), .ZN(n607) );
  INV_X2 U4346 ( .A(n608), .ZN(n981) );
  INV_X2 U4347 ( .A(n602), .ZN(n600) );
  INV_X2 U4348 ( .A(n601), .ZN(n980) );
  INV_X2 U4349 ( .A(n3640), .ZN(n3292) );
  INV_X2 U4350 ( .A(n333), .ZN(n3288) );
  INV_X2 U4351 ( .A(n3681), .ZN(n3287) );
  INV_X2 U4352 ( .A(n3603), .ZN(n3285) );
  INV_X2 U4353 ( .A(n3571), .ZN(n3284) );
  INV_X2 U4354 ( .A(n354), .ZN(n3281) );
  INV_X2 U4355 ( .A(n357), .ZN(n3280) );
  NAND2_X2 U4356 ( .A1(n3640), .A2(n3444), .ZN(n3195) );
  NAND2_X2 U4357 ( .A1(n3425), .A2(n3444), .ZN(n3162) );
  NAND2_X2 U4358 ( .A1(n327), .A2(n3444), .ZN(n3129) );
  NAND2_X2 U4359 ( .A1(n3795), .A2(n3444), .ZN(n3096) );
  NAND2_X2 U4360 ( .A1(n333), .A2(n3444), .ZN(n3063) );
  NAND2_X2 U4361 ( .A1(n3681), .A2(n3444), .ZN(n3030) );
  NAND2_X2 U4362 ( .A1(n339), .A2(n3444), .ZN(n2997) );
  NAND2_X2 U4363 ( .A1(n3603), .A2(n3444), .ZN(n2964) );
  NAND2_X2 U4364 ( .A1(n3571), .A2(n3444), .ZN(n2931) );
  NAND2_X2 U4365 ( .A1(n348), .A2(n3444), .ZN(n2898) );
  NAND2_X2 U4366 ( .A1(n3775), .A2(n3444), .ZN(n2865) );
  NAND2_X2 U4367 ( .A1(n354), .A2(n3444), .ZN(n2832) );
  NAND2_X2 U4368 ( .A1(n360), .A2(n3444), .ZN(n2766) );
  NAND2_X2 U4369 ( .A1(n363), .A2(n3444), .ZN(n2733) );
  NAND2_X2 U4370 ( .A1(n366), .A2(n3444), .ZN(n2700) );
  NOR2_X2 U4371 ( .A1(n3573), .A2(n3444), .ZN(n2603) );
  NOR2_X2 U4372 ( .A1(n3674), .A2(n3444), .ZN(n2569) );
  NOR2_X2 U4373 ( .A1(n3679), .A2(n3444), .ZN(n2535) );
  NOR2_X2 U4374 ( .A1(n3657), .A2(n3444), .ZN(n2501) );
  NOR2_X2 U4375 ( .A1(n3736), .A2(n3444), .ZN(n2433) );
  NOR2_X2 U4376 ( .A1(n3625), .A2(n3444), .ZN(n2399) );
  NOR2_X2 U4377 ( .A1(n393), .A2(n3444), .ZN(n2365) );
  NOR2_X2 U4378 ( .A1(n3728), .A2(n3444), .ZN(n2331) );
  NOR2_X2 U4379 ( .A1(n3613), .A2(n3444), .ZN(n2297) );
  NOR2_X2 U4380 ( .A1(n402), .A2(n3444), .ZN(n2263) );
  NOR2_X2 U4381 ( .A1(n3581), .A2(n3444), .ZN(n2229) );
  NOR2_X2 U4382 ( .A1(n3741), .A2(n3444), .ZN(n2195) );
  NOR2_X2 U4383 ( .A1(n3545), .A2(n3444), .ZN(n2161) );
  INV_X2 U4384 ( .A(n1486), .ZN(n1487) );
  INV_X2 U4385 ( .A(n1428), .ZN(n1429) );
  INV_X2 U4386 ( .A(n1374), .ZN(n1375) );
  INV_X2 U4387 ( .A(n1324), .ZN(n1325) );
  INV_X2 U4388 ( .A(n1278), .ZN(n1279) );
  INV_X2 U4389 ( .A(n1236), .ZN(n1237) );
  INV_X2 U4390 ( .A(n1198), .ZN(n1199) );
  INV_X2 U4391 ( .A(n1164), .ZN(n1165) );
  INV_X2 U4392 ( .A(n1134), .ZN(n1135) );
  INV_X2 U4393 ( .A(n1108), .ZN(n1109) );
  INV_X2 U4394 ( .A(n1086), .ZN(n1087) );
  INV_X2 U4395 ( .A(n1068), .ZN(n1069) );
  INV_X2 U4396 ( .A(n1054), .ZN(n1055) );
  INV_X2 U4397 ( .A(n1044), .ZN(n1045) );
  XOR2_X1 U4398 ( .A(n3817), .B(n3818), .Z(n1041) );
  XOR2_X1 U4399 ( .A(n2077), .B(n1044), .Z(n3818) );
  INV_X2 U4400 ( .A(n977), .ZN(n1040) );
  INV_X2 U4401 ( .A(n974), .ZN(n972) );
  INV_X2 U4402 ( .A(n969), .ZN(n1038) );
  INV_X2 U4403 ( .A(n966), .ZN(n964) );
  INV_X2 U4404 ( .A(n961), .ZN(n1036) );
  INV_X2 U4405 ( .A(n958), .ZN(n956) );
  INV_X2 U4406 ( .A(n952), .ZN(n950) );
  INV_X2 U4407 ( .A(n947), .ZN(n945) );
  INV_X2 U4408 ( .A(n940), .ZN(n938) );
  INV_X2 U4409 ( .A(n934), .ZN(n932) );
  INV_X2 U4410 ( .A(n929), .ZN(n927) );
  INV_X2 U4411 ( .A(n921), .ZN(n1029) );
  INV_X2 U4412 ( .A(n918), .ZN(n1028) );
  INV_X2 U4413 ( .A(n912), .ZN(n910) );
  INV_X2 U4414 ( .A(n907), .ZN(n1026) );
  INV_X2 U4415 ( .A(n902), .ZN(n900) );
  INV_X2 U4416 ( .A(n890), .ZN(n892) );
  INV_X2 U4417 ( .A(n880), .ZN(n1022) );
  INV_X2 U4418 ( .A(n874), .ZN(n872) );
  INV_X2 U4419 ( .A(n869), .ZN(n1020) );
  INV_X2 U4420 ( .A(n864), .ZN(n1019) );
  INV_X2 U4421 ( .A(n849), .ZN(n851) );
  INV_X2 U4422 ( .A(n846), .ZN(n844) );
  INV_X2 U4423 ( .A(n824), .ZN(n822) );
  INV_X2 U4424 ( .A(n3782), .ZN(n1002) );
  INV_X2 U4425 ( .A(n759), .ZN(n757) );
endmodule


module mul32_0_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n321, n324, n327, n330, n333, n336, n339, n342, n345, n348, n351,
         n354, n357, n360, n363, n366, n369, n372, n375, n381, n387, n390,
         n393, n396, n399, n405, n411, n414, n416, n419, n422, n425, n428,
         n431, n434, n440, n443, n446, n449, n455, n458, n461, n464, n465,
         n469, n471, n473, n475, n477, n479, n481, n483, n485, n487, n489,
         n491, n493, n495, n497, n499, n501, n503, n505, n507, n509, n511,
         n513, n515, n517, n519, n521, n523, n525, n527, n529, n531, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n600,
         n601, n602, n603, n604, n605, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n620, n621, n622, n623, n624,
         n625, n627, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n667, n668, n669, n670, n671, n672, n673,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n714, n715, n716, n717, n718, n719, n721, n724,
         n725, n726, n728, n729, n730, n731, n732, n734, n735, n736, n737,
         n738, n739, n744, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1003, n1004, n1005, n1006, n1008, n1009, n1010, n1011, n1012, n1018,
         n1019, n1020, n1022, n1026, n1028, n1029, n1036, n1038, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3228, n3229, n3230, n3232, n3233, n3234, n3235, n3236,
         n3240, n3241, n3242, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3290, n3291, n3292, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788;
  assign n321 = a[1];
  assign n324 = a[3];
  assign n327 = a[5];
  assign n330 = a[7];
  assign n333 = a[9];
  assign n336 = a[11];
  assign n339 = a[13];
  assign n342 = a[15];
  assign n345 = a[17];
  assign n348 = a[19];
  assign n351 = a[21];
  assign n354 = a[23];
  assign n357 = a[25];
  assign n360 = a[27];
  assign n363 = a[29];
  assign n366 = a[31];
  assign n465 = b[0];
  assign n469 = b[1];
  assign n471 = b[2];
  assign n473 = b[3];
  assign n475 = b[4];
  assign n477 = b[5];
  assign n479 = b[6];
  assign n481 = b[7];
  assign n483 = b[8];
  assign n485 = b[9];
  assign n487 = b[10];
  assign n489 = b[11];
  assign n491 = b[12];
  assign n493 = b[13];
  assign n495 = b[14];
  assign n497 = b[15];
  assign n499 = b[16];
  assign n501 = b[17];
  assign n503 = b[18];
  assign n505 = b[19];
  assign n507 = b[20];
  assign n509 = b[21];
  assign n511 = b[22];
  assign n513 = b[23];
  assign n515 = b[24];
  assign n517 = b[25];
  assign n519 = b[26];
  assign n521 = b[27];
  assign n523 = b[28];
  assign n525 = b[29];
  assign n527 = b[30];
  assign n529 = b[31];

  NAND2_X4 U322 ( .A1(n979), .A2(n597), .ZN(n533) );
  NOR2_X4 U324 ( .A1(n1043), .A2(n1046), .ZN(n596) );
  NAND2_X4 U325 ( .A1(n1043), .A2(n1046), .ZN(n597) );
  NAND2_X4 U330 ( .A1(n980), .A2(n602), .ZN(n534) );
  NOR2_X4 U332 ( .A1(n1050), .A2(n1047), .ZN(n601) );
  NAND2_X4 U333 ( .A1(n1050), .A2(n1047), .ZN(n602) );
  XOR2_X2 U334 ( .A(n610), .B(n535), .Z(product[60]) );
  NAND2_X4 U340 ( .A1(n981), .A2(n609), .ZN(n535) );
  NOR2_X4 U342 ( .A1(n1051), .A2(n1056), .ZN(n608) );
  NAND2_X4 U343 ( .A1(n1051), .A2(n1056), .ZN(n609) );
  NOR2_X4 U350 ( .A1(n633), .A2(n617), .ZN(n615) );
  NAND2_X4 U352 ( .A1(n983), .A2(n982), .ZN(n617) );
  AOI21_X4 U353 ( .B1(n982), .B2(n627), .A(n620), .ZN(n618) );
  NAND2_X4 U356 ( .A1(n982), .A2(n622), .ZN(n536) );
  NOR2_X4 U358 ( .A1(n1057), .A2(n1062), .ZN(n621) );
  NAND2_X4 U359 ( .A1(n1057), .A2(n1062), .ZN(n622) );
  NAND2_X4 U366 ( .A1(n983), .A2(n625), .ZN(n537) );
  NOR2_X4 U368 ( .A1(n1063), .A2(n1070), .ZN(n624) );
  NAND2_X4 U369 ( .A1(n1063), .A2(n1070), .ZN(n625) );
  NAND2_X4 U374 ( .A1(n673), .A2(n635), .ZN(n633) );
  NOR2_X4 U376 ( .A1(n656), .A2(n637), .ZN(n635) );
  NAND2_X4 U378 ( .A1(n646), .A2(n984), .ZN(n637) );
  AOI21_X4 U379 ( .B1(n647), .B2(n984), .A(n640), .ZN(n638) );
  NAND2_X4 U382 ( .A1(n984), .A2(n642), .ZN(n538) );
  NOR2_X4 U384 ( .A1(n1071), .A2(n1078), .ZN(n641) );
  NAND2_X4 U385 ( .A1(n1071), .A2(n1078), .ZN(n642) );
  NOR2_X4 U390 ( .A1(n651), .A2(n648), .ZN(n646) );
  OAI21_X4 U391 ( .B1(n648), .B2(n652), .A(n649), .ZN(n647) );
  NAND2_X4 U392 ( .A1(n985), .A2(n649), .ZN(n539) );
  NOR2_X4 U394 ( .A1(n1079), .A2(n1088), .ZN(n648) );
  NAND2_X4 U395 ( .A1(n1079), .A2(n1088), .ZN(n649) );
  NAND2_X4 U398 ( .A1(n986), .A2(n652), .ZN(n540) );
  NOR2_X4 U400 ( .A1(n1089), .A2(n1098), .ZN(n651) );
  NAND2_X4 U401 ( .A1(n1089), .A2(n1098), .ZN(n652) );
  NAND2_X4 U406 ( .A1(n658), .A2(n989), .ZN(n656) );
  NOR2_X4 U408 ( .A1(n663), .A2(n660), .ZN(n658) );
  OAI21_X4 U409 ( .B1(n660), .B2(n664), .A(n661), .ZN(n659) );
  NAND2_X4 U410 ( .A1(n987), .A2(n661), .ZN(n541) );
  NOR2_X4 U412 ( .A1(n1099), .A2(n1110), .ZN(n660) );
  NAND2_X4 U413 ( .A1(n1099), .A2(n1110), .ZN(n661) );
  NAND2_X4 U416 ( .A1(n988), .A2(n664), .ZN(n542) );
  NOR2_X4 U418 ( .A1(n1111), .A2(n1122), .ZN(n663) );
  NAND2_X4 U419 ( .A1(n1111), .A2(n1122), .ZN(n664) );
  NAND2_X4 U424 ( .A1(n989), .A2(n669), .ZN(n543) );
  NOR2_X4 U434 ( .A1(n680), .A2(n677), .ZN(n673) );
  OAI21_X4 U435 ( .B1(n677), .B2(n681), .A(n678), .ZN(n676) );
  NAND2_X4 U436 ( .A1(n990), .A2(n678), .ZN(n544) );
  NOR2_X4 U438 ( .A1(n1137), .A2(n1150), .ZN(n677) );
  NAND2_X4 U439 ( .A1(n1137), .A2(n1150), .ZN(n678) );
  NAND2_X4 U442 ( .A1(n991), .A2(n681), .ZN(n545) );
  NOR2_X4 U444 ( .A1(n1151), .A2(n1166), .ZN(n680) );
  NAND2_X4 U445 ( .A1(n1151), .A2(n1166), .ZN(n681) );
  NOR2_X4 U455 ( .A1(n692), .A2(n711), .ZN(n690) );
  AOI21_X4 U458 ( .B1(n694), .B2(n703), .A(n695), .ZN(n693) );
  NOR2_X4 U459 ( .A1(n699), .A2(n696), .ZN(n694) );
  OAI21_X4 U460 ( .B1(n696), .B2(n700), .A(n697), .ZN(n695) );
  NAND2_X4 U461 ( .A1(n992), .A2(n697), .ZN(n546) );
  NOR2_X4 U463 ( .A1(n1167), .A2(n1182), .ZN(n696) );
  NAND2_X4 U464 ( .A1(n1167), .A2(n1182), .ZN(n697) );
  NAND2_X4 U467 ( .A1(n993), .A2(n700), .ZN(n547) );
  NOR2_X4 U469 ( .A1(n1183), .A2(n1200), .ZN(n699) );
  NAND2_X4 U470 ( .A1(n1183), .A2(n1200), .ZN(n700) );
  NOR2_X4 U477 ( .A1(n1201), .A2(n1218), .ZN(n704) );
  NAND2_X4 U478 ( .A1(n1201), .A2(n1218), .ZN(n705) );
  NAND2_X4 U481 ( .A1(n725), .A2(n709), .ZN(n707) );
  NAND2_X4 U499 ( .A1(n996), .A2(n719), .ZN(n550) );
  NOR2_X4 U501 ( .A1(n1239), .A2(n1258), .ZN(n718) );
  NAND2_X4 U502 ( .A1(n1239), .A2(n1258), .ZN(n719) );
  NAND2_X4 U515 ( .A1(n997), .A2(n3654), .ZN(n551) );
  NAND2_X4 U533 ( .A1(n999), .A2(n748), .ZN(n553) );
  XOR2_X2 U537 ( .A(n756), .B(n554), .Z(product[41]) );
  NAND2_X4 U551 ( .A1(n757), .A2(n760), .ZN(n555) );
  XOR2_X2 U582 ( .A(n782), .B(n559), .Z(product[36]) );
  XNOR2_X2 U599 ( .A(n795), .B(n561), .ZN(product[34]) );
  AOI21_X4 U600 ( .B1(n795), .B2(n791), .A(n792), .ZN(n790) );
  XNOR2_X2 U607 ( .A(n802), .B(n562), .ZN(product[33]) );
  OAI21_X4 U608 ( .B1(n805), .B2(n796), .A(n797), .ZN(n795) );
  NAND2_X4 U613 ( .A1(n1008), .A2(n801), .ZN(n562) );
  XOR2_X2 U617 ( .A(n805), .B(n563), .Z(product[32]) );
  XNOR2_X2 U623 ( .A(n813), .B(n564), .ZN(product[31]) );
  NAND2_X4 U630 ( .A1(n1010), .A2(n812), .ZN(n564) );
  XOR2_X2 U634 ( .A(n816), .B(n565), .Z(product[30]) );
  XOR2_X2 U640 ( .A(n821), .B(n566), .Z(product[29]) );
  NAND2_X4 U644 ( .A1(n1012), .A2(n820), .ZN(n566) );
  XNOR2_X2 U648 ( .A(n826), .B(n567), .ZN(product[28]) );
  AOI21_X4 U649 ( .B1(n826), .B2(n822), .A(n823), .ZN(n821) );
  NAND2_X4 U652 ( .A1(n822), .A2(n825), .ZN(n567) );
  XOR2_X2 U656 ( .A(n836), .B(n568), .Z(product[27]) );
  NAND2_X4 U665 ( .A1(n832), .A2(n835), .ZN(n568) );
  XNOR2_X2 U669 ( .A(n841), .B(n569), .ZN(product[26]) );
  NAND2_X4 U673 ( .A1(n837), .A2(n840), .ZN(n569) );
  XNOR2_X2 U677 ( .A(n848), .B(n570), .ZN(product[25]) );
  XOR2_X2 U687 ( .A(n855), .B(n571), .Z(product[24]) );
  XNOR2_X2 U697 ( .A(n863), .B(n572), .ZN(product[23]) );
  NAND2_X4 U704 ( .A1(n1018), .A2(n862), .ZN(n572) );
  XOR2_X2 U708 ( .A(n866), .B(n573), .Z(product[22]) );
  NAND2_X4 U710 ( .A1(n1019), .A2(n865), .ZN(n573) );
  XOR2_X2 U714 ( .A(n871), .B(n574), .Z(product[21]) );
  AOI21_X4 U715 ( .B1(n876), .B2(n867), .A(n868), .ZN(n866) );
  NOR2_X4 U716 ( .A1(n869), .A2(n874), .ZN(n867) );
  OAI21_X4 U717 ( .B1(n869), .B2(n875), .A(n870), .ZN(n868) );
  NAND2_X4 U718 ( .A1(n1020), .A2(n870), .ZN(n574) );
  NOR2_X4 U720 ( .A1(n1862), .A2(n1881), .ZN(n869) );
  XNOR2_X2 U722 ( .A(n876), .B(n575), .ZN(product[20]) );
  AOI21_X4 U723 ( .B1(n876), .B2(n872), .A(n873), .ZN(n871) );
  NAND2_X4 U726 ( .A1(n872), .A2(n875), .ZN(n575) );
  NOR2_X4 U728 ( .A1(n1882), .A2(n1899), .ZN(n874) );
  NAND2_X4 U729 ( .A1(n1882), .A2(n1899), .ZN(n875) );
  XNOR2_X2 U730 ( .A(n882), .B(n576), .ZN(product[19]) );
  NOR2_X4 U733 ( .A1(n883), .A2(n880), .ZN(n878) );
  NAND2_X4 U735 ( .A1(n1022), .A2(n881), .ZN(n576) );
  NOR2_X4 U737 ( .A1(n1900), .A2(n1917), .ZN(n880) );
  NAND2_X4 U738 ( .A1(n1900), .A2(n1917), .ZN(n881) );
  XNOR2_X2 U739 ( .A(n889), .B(n577), .ZN(product[18]) );
  NAND2_X4 U741 ( .A1(n885), .A2(n892), .ZN(n883) );
  NAND2_X4 U745 ( .A1(n885), .A2(n888), .ZN(n577) );
  XOR2_X2 U749 ( .A(n896), .B(n578), .Z(product[17]) );
  OAI21_X4 U750 ( .B1(n896), .B2(n890), .A(n891), .ZN(n889) );
  NAND2_X4 U755 ( .A1(n892), .A2(n891), .ZN(n578) );
  NOR2_X4 U757 ( .A1(n1934), .A2(n1949), .ZN(n890) );
  NAND2_X4 U758 ( .A1(n1934), .A2(n1949), .ZN(n891) );
  XOR2_X2 U759 ( .A(n904), .B(n579), .Z(product[16]) );
  NAND2_X4 U766 ( .A1(n900), .A2(n903), .ZN(n579) );
  NOR2_X4 U768 ( .A1(n1950), .A2(n1963), .ZN(n902) );
  NAND2_X4 U769 ( .A1(n1950), .A2(n1963), .ZN(n903) );
  XOR2_X2 U770 ( .A(n909), .B(n580), .Z(product[15]) );
  AOI21_X4 U771 ( .B1(n914), .B2(n905), .A(n906), .ZN(n904) );
  NOR2_X4 U772 ( .A1(n907), .A2(n912), .ZN(n905) );
  OAI21_X4 U773 ( .B1(n907), .B2(n913), .A(n908), .ZN(n906) );
  NAND2_X4 U774 ( .A1(n1026), .A2(n908), .ZN(n580) );
  NOR2_X4 U776 ( .A1(n1964), .A2(n1977), .ZN(n907) );
  NAND2_X4 U777 ( .A1(n1964), .A2(n1977), .ZN(n908) );
  XNOR2_X2 U778 ( .A(n914), .B(n581), .ZN(product[14]) );
  AOI21_X4 U779 ( .B1(n914), .B2(n910), .A(n911), .ZN(n909) );
  NAND2_X4 U782 ( .A1(n910), .A2(n913), .ZN(n581) );
  NOR2_X4 U784 ( .A1(n1978), .A2(n1989), .ZN(n912) );
  NAND2_X4 U785 ( .A1(n1978), .A2(n1989), .ZN(n913) );
  XNOR2_X2 U786 ( .A(n920), .B(n582), .ZN(product[13]) );
  AOI21_X4 U788 ( .B1(n916), .B2(n924), .A(n917), .ZN(n915) );
  NOR2_X4 U789 ( .A1(n918), .A2(n921), .ZN(n916) );
  OAI21_X4 U790 ( .B1(n918), .B2(n922), .A(n919), .ZN(n917) );
  NAND2_X4 U791 ( .A1(n1028), .A2(n919), .ZN(n582) );
  NOR2_X4 U793 ( .A1(n1990), .A2(n2001), .ZN(n918) );
  NAND2_X4 U794 ( .A1(n1990), .A2(n2001), .ZN(n919) );
  XOR2_X2 U795 ( .A(n923), .B(n583), .Z(product[12]) );
  OAI21_X4 U796 ( .B1(n923), .B2(n921), .A(n922), .ZN(n920) );
  NAND2_X4 U797 ( .A1(n1029), .A2(n922), .ZN(n583) );
  NOR2_X4 U799 ( .A1(n2002), .A2(n2011), .ZN(n921) );
  NAND2_X4 U800 ( .A1(n2002), .A2(n2011), .ZN(n922) );
  XOR2_X2 U801 ( .A(n931), .B(n584), .Z(product[11]) );
  OAI21_X4 U803 ( .B1(n925), .B2(n937), .A(n926), .ZN(n924) );
  NAND2_X4 U804 ( .A1(n932), .A2(n927), .ZN(n925) );
  AOI21_X4 U805 ( .B1(n927), .B2(n933), .A(n928), .ZN(n926) );
  NAND2_X4 U808 ( .A1(n927), .A2(n930), .ZN(n584) );
  NOR2_X4 U810 ( .A1(n2012), .A2(n2021), .ZN(n929) );
  NAND2_X4 U811 ( .A1(n2012), .A2(n2021), .ZN(n930) );
  XNOR2_X2 U812 ( .A(n585), .B(n936), .ZN(product[10]) );
  AOI21_X4 U813 ( .B1(n936), .B2(n932), .A(n933), .ZN(n931) );
  NAND2_X4 U816 ( .A1(n932), .A2(n935), .ZN(n585) );
  NOR2_X4 U818 ( .A1(n2022), .A2(n2029), .ZN(n934) );
  NAND2_X4 U819 ( .A1(n2022), .A2(n2029), .ZN(n935) );
  XNOR2_X2 U820 ( .A(n586), .B(n942), .ZN(product[9]) );
  AOI21_X4 U822 ( .B1(n942), .B2(n938), .A(n939), .ZN(n937) );
  NAND2_X4 U825 ( .A1(n938), .A2(n941), .ZN(n586) );
  NOR2_X4 U827 ( .A1(n2030), .A2(n2037), .ZN(n940) );
  NAND2_X4 U828 ( .A1(n2030), .A2(n2037), .ZN(n941) );
  XOR2_X2 U829 ( .A(n949), .B(n587), .Z(product[8]) );
  OAI21_X4 U830 ( .B1(n943), .B2(n955), .A(n944), .ZN(n942) );
  NAND2_X4 U831 ( .A1(n945), .A2(n950), .ZN(n943) );
  AOI21_X4 U832 ( .B1(n945), .B2(n951), .A(n946), .ZN(n944) );
  NAND2_X4 U835 ( .A1(n945), .A2(n948), .ZN(n587) );
  NOR2_X4 U837 ( .A1(n2038), .A2(n2043), .ZN(n947) );
  NAND2_X4 U838 ( .A1(n2038), .A2(n2043), .ZN(n948) );
  XNOR2_X2 U839 ( .A(n954), .B(n588), .ZN(product[7]) );
  AOI21_X4 U840 ( .B1(n954), .B2(n950), .A(n951), .ZN(n949) );
  NAND2_X4 U843 ( .A1(n950), .A2(n953), .ZN(n588) );
  NOR2_X4 U845 ( .A1(n2044), .A2(n2049), .ZN(n952) );
  NAND2_X4 U846 ( .A1(n2044), .A2(n2049), .ZN(n953) );
  XNOR2_X2 U847 ( .A(n589), .B(n960), .ZN(product[6]) );
  AOI21_X4 U849 ( .B1(n956), .B2(n960), .A(n957), .ZN(n955) );
  NAND2_X4 U852 ( .A1(n956), .A2(n959), .ZN(n589) );
  NOR2_X4 U854 ( .A1(n2050), .A2(n2053), .ZN(n958) );
  NAND2_X4 U855 ( .A1(n2050), .A2(n2053), .ZN(n959) );
  XOR2_X2 U856 ( .A(n590), .B(n963), .Z(product[5]) );
  OAI21_X4 U857 ( .B1(n961), .B2(n963), .A(n962), .ZN(n960) );
  NAND2_X4 U858 ( .A1(n1036), .A2(n962), .ZN(n590) );
  NOR2_X4 U860 ( .A1(n2054), .A2(n2057), .ZN(n961) );
  NAND2_X4 U861 ( .A1(n2054), .A2(n2057), .ZN(n962) );
  XNOR2_X2 U862 ( .A(n591), .B(n968), .ZN(product[4]) );
  AOI21_X4 U863 ( .B1(n964), .B2(n968), .A(n965), .ZN(n963) );
  NAND2_X4 U866 ( .A1(n964), .A2(n967), .ZN(n591) );
  NOR2_X4 U868 ( .A1(n2058), .A2(n2059), .ZN(n966) );
  NAND2_X4 U869 ( .A1(n2058), .A2(n2059), .ZN(n967) );
  XOR2_X2 U870 ( .A(n592), .B(n971), .Z(product[3]) );
  OAI21_X4 U871 ( .B1(n969), .B2(n971), .A(n970), .ZN(n968) );
  NAND2_X4 U872 ( .A1(n1038), .A2(n970), .ZN(n592) );
  NOR2_X4 U874 ( .A1(n2060), .A2(n2075), .ZN(n969) );
  NAND2_X4 U875 ( .A1(n2060), .A2(n2075), .ZN(n970) );
  XNOR2_X2 U876 ( .A(n593), .B(n976), .ZN(product[2]) );
  AOI21_X4 U877 ( .B1(n972), .B2(n976), .A(n973), .ZN(n971) );
  NAND2_X4 U880 ( .A1(n972), .A2(n975), .ZN(n593) );
  NOR2_X4 U882 ( .A1(n2603), .A2(n2635), .ZN(n974) );
  NAND2_X4 U883 ( .A1(n2603), .A2(n2635), .ZN(n975) );
  NAND2_X4 U886 ( .A1(n1040), .A2(n978), .ZN(n594) );
  NOR2_X4 U888 ( .A1(n2636), .A2(n2076), .ZN(n977) );
  NAND2_X4 U889 ( .A1(n2636), .A2(n2076), .ZN(n978) );
  FA_X1 U890 ( .A(n2095), .B(n1045), .CI(n1048), .CO(n1042), .S(n1043) );
  FA_X1 U892 ( .A(n1052), .B(n2128), .CI(n1049), .CO(n1046), .S(n1047) );
  FA_X1 U893 ( .A(n2078), .B(n1054), .CI(n2096), .CO(n1048), .S(n1049) );
  FA_X1 U894 ( .A(n1053), .B(n1060), .CI(n1058), .CO(n1050), .S(n1051) );
  FA_X1 U895 ( .A(n2129), .B(n1055), .CI(n2097), .CO(n1052), .S(n1053) );
  FA_X1 U897 ( .A(n1064), .B(n1061), .CI(n1059), .CO(n1056), .S(n1057) );
  FA_X1 U898 ( .A(n2162), .B(n2098), .CI(n1066), .CO(n1058), .S(n1059) );
  FA_X1 U899 ( .A(n2079), .B(n1068), .CI(n2130), .CO(n1060), .S(n1061) );
  FA_X1 U900 ( .A(n1072), .B(n1067), .CI(n1065), .CO(n1062), .S(n1063) );
  FA_X1 U901 ( .A(n1076), .B(n2099), .CI(n1074), .CO(n1064), .S(n1065) );
  FA_X1 U902 ( .A(n2163), .B(n1069), .CI(n2131), .CO(n1066), .S(n1067) );
  FA_X1 U904 ( .A(n1080), .B(n1082), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U905 ( .A(n1077), .B(n1084), .CI(n1075), .CO(n1072), .S(n1073) );
  FA_X1 U906 ( .A(n2132), .B(n2100), .CI(n2196), .CO(n1074), .S(n1075) );
  FA_X1 U907 ( .A(n2080), .B(n1086), .CI(n2164), .CO(n1076), .S(n1077) );
  FA_X1 U908 ( .A(n1090), .B(n1083), .CI(n1081), .CO(n1078), .S(n1079) );
  FA_X1 U909 ( .A(n1085), .B(n1094), .CI(n1092), .CO(n1080), .S(n1081) );
  FA_X1 U910 ( .A(n2101), .B(n2133), .CI(n1096), .CO(n1082), .S(n1083) );
  FA_X1 U911 ( .A(n2197), .B(n1087), .CI(n2165), .CO(n1084), .S(n1085) );
  FA_X1 U913 ( .A(n1100), .B(n1093), .CI(n1091), .CO(n1088), .S(n1089) );
  FA_X1 U914 ( .A(n1095), .B(n1097), .CI(n1102), .CO(n1090), .S(n1091) );
  FA_X1 U915 ( .A(n1106), .B(n2230), .CI(n1104), .CO(n1092), .S(n1093) );
  FA_X1 U916 ( .A(n2102), .B(n2134), .CI(n2198), .CO(n1094), .S(n1095) );
  FA_X1 U917 ( .A(n2081), .B(n1108), .CI(n2166), .CO(n1096), .S(n1097) );
  FA_X1 U918 ( .A(n1112), .B(n1103), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U919 ( .A(n1116), .B(n1105), .CI(n1114), .CO(n1100), .S(n1101) );
  FA_X1 U920 ( .A(n1118), .B(n1120), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U921 ( .A(n2135), .B(n2103), .CI(n2167), .CO(n1104), .S(n1105) );
  FA_X1 U922 ( .A(n2231), .B(n1109), .CI(n2199), .CO(n1106), .S(n1107) );
  FA_X1 U924 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U925 ( .A(n1117), .B(n1128), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U926 ( .A(n1121), .B(n1130), .CI(n1119), .CO(n1114), .S(n1115) );
  FA_X1 U927 ( .A(n2264), .B(n2136), .CI(n1132), .CO(n1116), .S(n1117) );
  FA_X1 U928 ( .A(n2104), .B(n2168), .CI(n2232), .CO(n1118), .S(n1119) );
  FA_X1 U929 ( .A(n2082), .B(n1134), .CI(n2200), .CO(n1120), .S(n1121) );
  FA_X1 U930 ( .A(n1138), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U931 ( .A(n1129), .B(n1142), .CI(n1140), .CO(n1124), .S(n1125) );
  FA_X1 U932 ( .A(n1133), .B(n1144), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U933 ( .A(n1148), .B(n2137), .CI(n1146), .CO(n1128), .S(n1129) );
  FA_X1 U934 ( .A(n2105), .B(n2201), .CI(n2169), .CO(n1130), .S(n1131) );
  FA_X1 U935 ( .A(n2265), .B(n1135), .CI(n2233), .CO(n1132), .S(n1133) );
  FA_X1 U937 ( .A(n1152), .B(n1141), .CI(n1139), .CO(n1136), .S(n1137) );
  FA_X1 U938 ( .A(n1143), .B(n1156), .CI(n1154), .CO(n1138), .S(n1139) );
  FA_X1 U939 ( .A(n1145), .B(n1147), .CI(n1158), .CO(n1140), .S(n1141) );
  FA_X1 U940 ( .A(n1160), .B(n1162), .CI(n1149), .CO(n1142), .S(n1143) );
  FA_X1 U941 ( .A(n2266), .B(n2106), .CI(n2298), .CO(n1144), .S(n1145) );
  FA_X1 U942 ( .A(n2138), .B(n2170), .CI(n2234), .CO(n1146), .S(n1147) );
  FA_X1 U943 ( .A(n2083), .B(n1164), .CI(n2202), .CO(n1148), .S(n1149) );
  FA_X1 U944 ( .A(n1168), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U945 ( .A(n1157), .B(n1172), .CI(n1170), .CO(n1152), .S(n1153) );
  FA_X1 U946 ( .A(n1174), .B(n1161), .CI(n1159), .CO(n1154), .S(n1155) );
  FA_X1 U947 ( .A(n1176), .B(n1178), .CI(n1163), .CO(n1156), .S(n1157) );
  FA_X1 U948 ( .A(n2171), .B(n2203), .CI(n1180), .CO(n1158), .S(n1159) );
  FA_X1 U949 ( .A(n2107), .B(n2235), .CI(n2139), .CO(n1160), .S(n1161) );
  FA_X1 U950 ( .A(n2299), .B(n1165), .CI(n2267), .CO(n1162), .S(n1163) );
  FA_X1 U952 ( .A(n1184), .B(n1171), .CI(n1169), .CO(n1166), .S(n1167) );
  FA_X1 U953 ( .A(n1173), .B(n1188), .CI(n1186), .CO(n1168), .S(n1169) );
  FA_X1 U954 ( .A(n1190), .B(n1179), .CI(n1175), .CO(n1170), .S(n1171) );
  FA_X1 U955 ( .A(n1181), .B(n1192), .CI(n1177), .CO(n1172), .S(n1173) );
  FA_X1 U956 ( .A(n1196), .B(n2332), .CI(n1194), .CO(n1174), .S(n1175) );
  FA_X1 U957 ( .A(n2268), .B(n2140), .CI(n2300), .CO(n1176), .S(n1177) );
  FA_X1 U958 ( .A(n2108), .B(n2204), .CI(n2172), .CO(n1178), .S(n1179) );
  FA_X1 U959 ( .A(n2084), .B(n1198), .CI(n2236), .CO(n1180), .S(n1181) );
  FA_X1 U960 ( .A(n1202), .B(n1187), .CI(n1185), .CO(n1182), .S(n1183) );
  FA_X1 U961 ( .A(n1189), .B(n1206), .CI(n1204), .CO(n1184), .S(n1185) );
  FA_X1 U962 ( .A(n1208), .B(n1210), .CI(n1191), .CO(n1186), .S(n1187) );
  FA_X1 U963 ( .A(n1193), .B(n1197), .CI(n1195), .CO(n1188), .S(n1189) );
  FA_X1 U964 ( .A(n1214), .B(n1216), .CI(n1212), .CO(n1190), .S(n1191) );
  FA_X1 U965 ( .A(n2141), .B(n2205), .CI(n2173), .CO(n1192), .S(n1193) );
  FA_X1 U966 ( .A(n2109), .B(n2269), .CI(n2237), .CO(n1194), .S(n1195) );
  FA_X1 U967 ( .A(n2333), .B(n1199), .CI(n2301), .CO(n1196), .S(n1197) );
  FA_X1 U969 ( .A(n1220), .B(n1205), .CI(n1203), .CO(n1200), .S(n1201) );
  FA_X1 U970 ( .A(n1207), .B(n1224), .CI(n1222), .CO(n1202), .S(n1203) );
  FA_X1 U971 ( .A(n1211), .B(n1226), .CI(n1209), .CO(n1204), .S(n1205) );
  FA_X1 U972 ( .A(n1215), .B(n1213), .CI(n1228), .CO(n1206), .S(n1207) );
  FA_X1 U973 ( .A(n1230), .B(n1232), .CI(n1217), .CO(n1208), .S(n1209) );
  FA_X1 U974 ( .A(n2366), .B(n2334), .CI(n1234), .CO(n1210), .S(n1211) );
  FA_X1 U975 ( .A(n2302), .B(n2174), .CI(n2270), .CO(n1212), .S(n1213) );
  FA_X1 U976 ( .A(n2142), .B(n2206), .CI(n2110), .CO(n1214), .S(n1215) );
  FA_X1 U977 ( .A(n2085), .B(n1236), .CI(n2238), .CO(n1216), .S(n1217) );
  FA_X1 U978 ( .A(n1240), .B(n1223), .CI(n1221), .CO(n1218), .S(n1219) );
  FA_X1 U979 ( .A(n1225), .B(n1244), .CI(n1242), .CO(n1220), .S(n1221) );
  FA_X1 U980 ( .A(n1246), .B(n1229), .CI(n1227), .CO(n1222), .S(n1223) );
  FA_X1 U981 ( .A(n1233), .B(n1231), .CI(n1248), .CO(n1224), .S(n1225) );
  FA_X1 U982 ( .A(n1250), .B(n1252), .CI(n1235), .CO(n1226), .S(n1227) );
  FA_X1 U983 ( .A(n1256), .B(n2239), .CI(n1254), .CO(n1228), .S(n1229) );
  FA_X1 U984 ( .A(n2175), .B(n2271), .CI(n2207), .CO(n1230), .S(n1231) );
  FA_X1 U985 ( .A(n2111), .B(n2303), .CI(n2143), .CO(n1232), .S(n1233) );
  FA_X1 U986 ( .A(n2367), .B(n1237), .CI(n2335), .CO(n1234), .S(n1235) );
  FA_X1 U988 ( .A(n1260), .B(n1243), .CI(n1241), .CO(n1238), .S(n1239) );
  FA_X1 U989 ( .A(n1245), .B(n1264), .CI(n1262), .CO(n1240), .S(n1241) );
  FA_X1 U990 ( .A(n1249), .B(n1266), .CI(n1247), .CO(n1242), .S(n1243) );
  FA_X1 U991 ( .A(n1270), .B(n1251), .CI(n1268), .CO(n1244), .S(n1245) );
  FA_X1 U992 ( .A(n1253), .B(n1257), .CI(n1255), .CO(n1246), .S(n1247) );
  FA_X1 U993 ( .A(n1272), .B(n1276), .CI(n1274), .CO(n1248), .S(n1249) );
  FA_X1 U994 ( .A(n2336), .B(n2368), .CI(n2400), .CO(n1250), .S(n1251) );
  FA_X1 U995 ( .A(n2304), .B(n2144), .CI(n2208), .CO(n1252), .S(n1253) );
  FA_X1 U996 ( .A(n2112), .B(n2240), .CI(n2176), .CO(n1254), .S(n1255) );
  FA_X1 U997 ( .A(n2086), .B(n1278), .CI(n2272), .CO(n1256), .S(n1257) );
  FA_X1 U998 ( .A(n1282), .B(n1263), .CI(n1261), .CO(n1258), .S(n1259) );
  FA_X1 U999 ( .A(n1265), .B(n1286), .CI(n1284), .CO(n1260), .S(n1261) );
  FA_X1 U1000 ( .A(n1269), .B(n1288), .CI(n1267), .CO(n1262), .S(n1263) );
  FA_X1 U1001 ( .A(n1271), .B(n1292), .CI(n1290), .CO(n1264), .S(n1265) );
  FA_X1 U1002 ( .A(n1273), .B(n1277), .CI(n1275), .CO(n1266), .S(n1267) );
  FA_X1 U1003 ( .A(n1294), .B(n1298), .CI(n1296), .CO(n1268), .S(n1269) );
  FA_X1 U1004 ( .A(n2273), .B(n2305), .CI(n1300), .CO(n1270), .S(n1271) );
  FA_X1 U1005 ( .A(n2177), .B(n2241), .CI(n2209), .CO(n1272), .S(n1273) );
  FA_X1 U1006 ( .A(n2113), .B(n2337), .CI(n2145), .CO(n1274), .S(n1275) );
  FA_X1 U1007 ( .A(n2401), .B(n1279), .CI(n2369), .CO(n1276), .S(n1277) );
  FA_X1 U1009 ( .A(n1285), .B(n1304), .CI(n1283), .CO(n1280), .S(n1281) );
  FA_X1 U1010 ( .A(n1287), .B(n1308), .CI(n1306), .CO(n1282), .S(n1283) );
  FA_X1 U1011 ( .A(n1310), .B(n1291), .CI(n1289), .CO(n1284), .S(n1285) );
  FA_X1 U1012 ( .A(n1312), .B(n1314), .CI(n1293), .CO(n1286), .S(n1287) );
  FA_X1 U1013 ( .A(n1299), .B(n1295), .CI(n1297), .CO(n1288), .S(n1289) );
  FA_X1 U1014 ( .A(n1316), .B(n1318), .CI(n1301), .CO(n1290), .S(n1291) );
  FA_X1 U1015 ( .A(n1322), .B(n2434), .CI(n1320), .CO(n1292), .S(n1293) );
  FA_X1 U1016 ( .A(n2210), .B(n2402), .CI(n2370), .CO(n1294), .S(n1295) );
  FA_X1 U1017 ( .A(n2178), .B(n2306), .CI(n2338), .CO(n1296), .S(n1297) );
  FA_X1 U1018 ( .A(n2114), .B(n2242), .CI(n2146), .CO(n1298), .S(n1299) );
  FA_X1 U1019 ( .A(n2087), .B(n1324), .CI(n2274), .CO(n1300), .S(n1301) );
  FA_X1 U1020 ( .A(n1328), .B(n1307), .CI(n1305), .CO(n1302), .S(n1303) );
  FA_X1 U1021 ( .A(n1309), .B(n1332), .CI(n1330), .CO(n1304), .S(n1305) );
  FA_X1 U1022 ( .A(n1334), .B(n1313), .CI(n1311), .CO(n1306), .S(n1307) );
  FA_X1 U1023 ( .A(n1315), .B(n1338), .CI(n1336), .CO(n1308), .S(n1309) );
  FA_X1 U1024 ( .A(n1321), .B(n1319), .CI(n1340), .CO(n1310), .S(n1311) );
  FA_X1 U1025 ( .A(n1323), .B(n1342), .CI(n1317), .CO(n1312), .S(n1313) );
  FA_X1 U1026 ( .A(n1346), .B(n1348), .CI(n1344), .CO(n1314), .S(n1315) );
  FA_X1 U1027 ( .A(n2243), .B(n2307), .CI(n2275), .CO(n1316), .S(n1317) );
  FA_X1 U1028 ( .A(n2339), .B(n2179), .CI(n2211), .CO(n1318), .S(n1319) );
  FA_X1 U1029 ( .A(n2115), .B(n2371), .CI(n2147), .CO(n1320), .S(n1321) );
  FA_X1 U1030 ( .A(n2435), .B(n1325), .CI(n2403), .CO(n1322), .S(n1323) );
  FA_X1 U1032 ( .A(n1352), .B(n1331), .CI(n1329), .CO(n1326), .S(n1327) );
  FA_X1 U1033 ( .A(n1333), .B(n1356), .CI(n1354), .CO(n1328), .S(n1329) );
  FA_X1 U1035 ( .A(n1360), .B(n1341), .CI(n1339), .CO(n1332), .S(n1333) );
  FA_X1 U1037 ( .A(n1343), .B(n1349), .CI(n1345), .CO(n1336), .S(n1337) );
  FA_X1 U1038 ( .A(n1366), .B(n1370), .CI(n1368), .CO(n1338), .S(n1339) );
  FA_X1 U1039 ( .A(n2468), .B(n2436), .CI(n1372), .CO(n1340), .S(n1341) );
  FA_X1 U1040 ( .A(n2212), .B(n2404), .CI(n2372), .CO(n1342), .S(n1343) );
  FA_X1 U1041 ( .A(n2116), .B(n2340), .CI(n2244), .CO(n1344), .S(n1345) );
  FA_X1 U1042 ( .A(n2148), .B(n2276), .CI(n2180), .CO(n1346), .S(n1347) );
  FA_X1 U1043 ( .A(n2088), .B(n1374), .CI(n2308), .CO(n1348), .S(n1349) );
  FA_X1 U1044 ( .A(n1378), .B(n1355), .CI(n1353), .CO(n1350), .S(n1351) );
  FA_X1 U1045 ( .A(n1357), .B(n1382), .CI(n1380), .CO(n1352), .S(n1353) );
  FA_X1 U1046 ( .A(n1384), .B(n1361), .CI(n1359), .CO(n1354), .S(n1355) );
  FA_X1 U1047 ( .A(n1386), .B(n1365), .CI(n1363), .CO(n1356), .S(n1357) );
  FA_X1 U1048 ( .A(n1390), .B(n1369), .CI(n1388), .CO(n1358), .S(n1359) );
  FA_X1 U1049 ( .A(n1367), .B(n1373), .CI(n1371), .CO(n1360), .S(n1361) );
  FA_X1 U1050 ( .A(n1394), .B(n1396), .CI(n1392), .CO(n1362), .S(n1363) );
  FA_X1 U1051 ( .A(n1400), .B(n2341), .CI(n1398), .CO(n1364), .S(n1365) );
  FA_X1 U1052 ( .A(n2245), .B(n2373), .CI(n2309), .CO(n1366), .S(n1367) );
  FA_X1 U1053 ( .A(n2181), .B(n2405), .CI(n2213), .CO(n1368), .S(n1369) );
  FA_X1 U1054 ( .A(n2117), .B(n2437), .CI(n2149), .CO(n1370), .S(n1371) );
  FA_X1 U1055 ( .A(n2469), .B(n1375), .CI(n2277), .CO(n1372), .S(n1373) );
  FA_X1 U1057 ( .A(n1404), .B(n1381), .CI(n1379), .CO(n1376), .S(n1377) );
  FA_X1 U1058 ( .A(n1383), .B(n1408), .CI(n1406), .CO(n1378), .S(n1379) );
  FA_X1 U1059 ( .A(n1410), .B(n1387), .CI(n1385), .CO(n1380), .S(n1381) );
  FA_X1 U1060 ( .A(n1389), .B(n1391), .CI(n1412), .CO(n1382), .S(n1383) );
  FA_X1 U1061 ( .A(n1416), .B(n1418), .CI(n1414), .CO(n1384), .S(n1385) );
  FA_X1 U1062 ( .A(n1399), .B(n1397), .CI(n1393), .CO(n1386), .S(n1387) );
  FA_X1 U1063 ( .A(n1401), .B(n1422), .CI(n1395), .CO(n1388), .S(n1389) );
  FA_X1 U1064 ( .A(n1420), .B(n1426), .CI(n1424), .CO(n1390), .S(n1391) );
  FA_X1 U1065 ( .A(n2438), .B(n2470), .CI(n2502), .CO(n1392), .S(n1393) );
  FA_X1 U1066 ( .A(n2406), .B(n2246), .CI(n2374), .CO(n1394), .S(n1395) );
  FA_X1 U1067 ( .A(n2118), .B(n2310), .CI(n2214), .CO(n1396), .S(n1397) );
  FA_X1 U1068 ( .A(n2182), .B(n2278), .CI(n2150), .CO(n1398), .S(n1399) );
  FA_X1 U1069 ( .A(n2089), .B(n1428), .CI(n2342), .CO(n1400), .S(n1401) );
  FA_X1 U1072 ( .A(n1438), .B(n1413), .CI(n1411), .CO(n1406), .S(n1407) );
  FA_X1 U1073 ( .A(n1415), .B(n1417), .CI(n1440), .CO(n1408), .S(n1409) );
  FA_X1 U1074 ( .A(n1419), .B(n1444), .CI(n1442), .CO(n1410), .S(n1411) );
  FA_X1 U1075 ( .A(n1425), .B(n1423), .CI(n1446), .CO(n1412), .S(n1413) );
  FA_X1 U1076 ( .A(n1427), .B(n1452), .CI(n1421), .CO(n1414), .S(n1415) );
  FA_X1 U1077 ( .A(n1448), .B(n1454), .CI(n1450), .CO(n1416), .S(n1417) );
  FA_X1 U1078 ( .A(n2247), .B(n2311), .CI(n1456), .CO(n1418), .S(n1419) );
  FA_X1 U1079 ( .A(n2183), .B(n2343), .CI(n2215), .CO(n1420), .S(n1421) );
  FA_X1 U1080 ( .A(n2375), .B(n2407), .CI(n2151), .CO(n1422), .S(n1423) );
  FA_X1 U1081 ( .A(n2439), .B(n2279), .CI(n2119), .CO(n1424), .S(n1425) );
  FA_X1 U1082 ( .A(n2503), .B(n1429), .CI(n2471), .CO(n1426), .S(n1427) );
  FA_X1 U1085 ( .A(n1437), .B(n1464), .CI(n1462), .CO(n1432), .S(n1433) );
  FA_X1 U1086 ( .A(n1466), .B(n1441), .CI(n1439), .CO(n1434), .S(n1435) );
  FA_X1 U1087 ( .A(n1443), .B(n1445), .CI(n1468), .CO(n1436), .S(n1437) );
  FA_X1 U1088 ( .A(n1472), .B(n1447), .CI(n1470), .CO(n1438), .S(n1439) );
  FA_X1 U1089 ( .A(n1453), .B(n1455), .CI(n1474), .CO(n1440), .S(n1441) );
  FA_X1 U1090 ( .A(n1449), .B(n1457), .CI(n1451), .CO(n1442), .S(n1443) );
  FA_X1 U1091 ( .A(n1482), .B(n1478), .CI(n1480), .CO(n1444), .S(n1445) );
  FA_X1 U1092 ( .A(n1484), .B(n2536), .CI(n1476), .CO(n1446), .S(n1447) );
  FA_X1 U1093 ( .A(n2504), .B(n2280), .CI(n2472), .CO(n1448), .S(n1449) );
  FA_X1 U1094 ( .A(n2248), .B(n2408), .CI(n2440), .CO(n1450), .S(n1451) );
  FA_X1 U1095 ( .A(n2152), .B(n2376), .CI(n2216), .CO(n1452), .S(n1453) );
  FA_X1 U1096 ( .A(n2120), .B(n2184), .CI(n2312), .CO(n1454), .S(n1455) );
  FA_X1 U1097 ( .A(n2090), .B(n1486), .CI(n2344), .CO(n1456), .S(n1457) );
  FA_X1 U1098 ( .A(n1490), .B(n1463), .CI(n1461), .CO(n1458), .S(n1459) );
  FA_X1 U1099 ( .A(n1465), .B(n1494), .CI(n1492), .CO(n1460), .S(n1461) );
  FA_X1 U1101 ( .A(n1471), .B(n1473), .CI(n1498), .CO(n1464), .S(n1465) );
  FA_X1 U1103 ( .A(n1506), .B(n1481), .CI(n1504), .CO(n1468), .S(n1469) );
  FA_X1 U1104 ( .A(n1483), .B(n1477), .CI(n1479), .CO(n1470), .S(n1471) );
  FA_X1 U1105 ( .A(n1514), .B(n1512), .CI(n1485), .CO(n1472), .S(n1473) );
  FA_X1 U1106 ( .A(n1508), .B(n1516), .CI(n1510), .CO(n1474), .S(n1475) );
  FA_X1 U1107 ( .A(n2313), .B(n2345), .CI(n2249), .CO(n1476), .S(n1477) );
  FA_X1 U1108 ( .A(n2185), .B(n2377), .CI(n2217), .CO(n1478), .S(n1479) );
  FA_X1 U1109 ( .A(n2153), .B(n2441), .CI(n2409), .CO(n1480), .S(n1481) );
  FA_X1 U1110 ( .A(n2473), .B(n2281), .CI(n2121), .CO(n1482), .S(n1483) );
  FA_X1 U1111 ( .A(n2537), .B(n1487), .CI(n2505), .CO(n1484), .S(n1485) );
  FA_X1 U1113 ( .A(n1493), .B(n1520), .CI(n1491), .CO(n1488), .S(n1489) );
  FA_X1 U1114 ( .A(n1522), .B(n1524), .CI(n1495), .CO(n1490), .S(n1491) );
  FA_X1 U1115 ( .A(n1499), .B(n1526), .CI(n1497), .CO(n1492), .S(n1493) );
  FA_X1 U1116 ( .A(n1501), .B(n1503), .CI(n1528), .CO(n1494), .S(n1495) );
  FA_X1 U1118 ( .A(n1534), .B(n1536), .CI(n1507), .CO(n1498), .S(n1499) );
  FA_X1 U1119 ( .A(n1515), .B(n1513), .CI(n1511), .CO(n1500), .S(n1501) );
  FA_X1 U1120 ( .A(n1517), .B(n1540), .CI(n1509), .CO(n1502), .S(n1503) );
  FA_X1 U1121 ( .A(n1544), .B(n1538), .CI(n1542), .CO(n1504), .S(n1505) );
  FA_X1 U1122 ( .A(n2570), .B(n2474), .CI(n1546), .CO(n1506), .S(n1507) );
  FA_X1 U1124 ( .A(n2346), .B(n2250), .CI(n2282), .CO(n1510), .S(n1511) );
  FA_X1 U1125 ( .A(n2218), .B(n2410), .CI(n2186), .CO(n1512), .S(n1513) );
  FA_X1 U1126 ( .A(n2154), .B(n2122), .CI(n2314), .CO(n1514), .S(n1515) );
  FA_X1 U1127 ( .A(n2091), .B(n1548), .CI(n2378), .CO(n1516), .S(n1517) );
  FA_X1 U1131 ( .A(n1531), .B(n1533), .CI(n1560), .CO(n1524), .S(n1525) );
  FA_X1 U1133 ( .A(n1566), .B(n1568), .CI(n1564), .CO(n1528), .S(n1529) );
  FA_X1 U1135 ( .A(n1547), .B(n1572), .CI(n1539), .CO(n1532), .S(n1533) );
  FA_X1 U1136 ( .A(n1576), .B(n1570), .CI(n1574), .CO(n1534), .S(n1535) );
  FA_X1 U1137 ( .A(n2411), .B(n2379), .CI(n1578), .CO(n1536), .S(n1537) );
  FA_X1 U1138 ( .A(n2315), .B(n2443), .CI(n2347), .CO(n1538), .S(n1539) );
  FA_X1 U1139 ( .A(n2475), .B(n2251), .CI(n2283), .CO(n1540), .S(n1541) );
  FA_X1 U1141 ( .A(n2123), .B(n2539), .CI(n2155), .CO(n1544), .S(n1545) );
  FA_X1 U1142 ( .A(n1580), .B(n2092), .CI(n2571), .CO(n1546), .S(n1547) );
  FA_X1 U1145 ( .A(n1557), .B(n1559), .CI(n1585), .CO(n1552), .S(n1553) );
  FA_X1 U1146 ( .A(n1561), .B(n1589), .CI(n1587), .CO(n1554), .S(n1555) );
  FA_X1 U1147 ( .A(n1591), .B(n1565), .CI(n1563), .CO(n1556), .S(n1557) );
  FA_X1 U1148 ( .A(n1593), .B(n1569), .CI(n1567), .CO(n1558), .S(n1559) );
  FA_X1 U1149 ( .A(n1597), .B(n1575), .CI(n1595), .CO(n1560), .S(n1561) );
  FA_X1 U1151 ( .A(n1599), .B(n1605), .CI(n1579), .CO(n1564), .S(n1565) );
  FA_X1 U1152 ( .A(n1607), .B(n1601), .CI(n1603), .CO(n1566), .S(n1567) );
  FA_X1 U1153 ( .A(n2604), .B(n2508), .CI(n1609), .CO(n1568), .S(n1569) );
  FA_X1 U1155 ( .A(n2284), .B(n2380), .CI(n2316), .CO(n1572), .S(n1573) );
  FA_X1 U1156 ( .A(n2220), .B(n2444), .CI(n2252), .CO(n1574), .S(n1575) );
  FA_X1 U1157 ( .A(n2188), .B(n2124), .CI(n2348), .CO(n1576), .S(n1577) );
  FA_X1 U1158 ( .A(n1580), .B(n2412), .CI(n2156), .CO(n1578), .S(n1579) );
  FA_X1 U1161 ( .A(n1588), .B(n1590), .CI(n1615), .CO(n1583), .S(n1584) );
  FA_X1 U1162 ( .A(n1619), .B(n1592), .CI(n1617), .CO(n1585), .S(n1586) );
  FA_X1 U1163 ( .A(n1621), .B(n1596), .CI(n1594), .CO(n1587), .S(n1588) );
  FA_X1 U1164 ( .A(n1623), .B(n1625), .CI(n1598), .CO(n1589), .S(n1590) );
  FA_X1 U1165 ( .A(n1600), .B(n1606), .CI(n1627), .CO(n1591), .S(n1592) );
  FA_X1 U1166 ( .A(n1604), .B(n1602), .CI(n1608), .CO(n1593), .S(n1594) );
  FA_X1 U1167 ( .A(n1633), .B(n1629), .CI(n1610), .CO(n1595), .S(n1596) );
  FA_X1 U1168 ( .A(n1637), .B(n1631), .CI(n1635), .CO(n1597), .S(n1598) );
  FA_X1 U1169 ( .A(n2445), .B(n2413), .CI(n1639), .CO(n1599), .S(n1600) );
  FA_X1 U1170 ( .A(n2349), .B(n2477), .CI(n2317), .CO(n1601), .S(n1602) );
  FA_X1 U1171 ( .A(n2285), .B(n2509), .CI(n2253), .CO(n1603), .S(n1604) );
  FA_X1 U1172 ( .A(n2541), .B(n2381), .CI(n2221), .CO(n1605), .S(n1606) );
  FA_X1 U1173 ( .A(n2189), .B(n2573), .CI(n2125), .CO(n1607), .S(n1608) );
  FA_X1 U1174 ( .A(n2157), .B(n2093), .CI(n2605), .CO(n1609), .S(n1610) );
  FA_X1 U1175 ( .A(n1643), .B(n1616), .CI(n1614), .CO(n1611), .S(n1612) );
  FA_X1 U1176 ( .A(n1618), .B(n1620), .CI(n1645), .CO(n1613), .S(n1614) );
  FA_X1 U1177 ( .A(n1649), .B(n1622), .CI(n1647), .CO(n1615), .S(n1616) );
  FA_X1 U1178 ( .A(n1651), .B(n1626), .CI(n1624), .CO(n1617), .S(n1618) );
  FA_X1 U1179 ( .A(n1628), .B(n1655), .CI(n1653), .CO(n1619), .S(n1620) );
  FA_X1 U1180 ( .A(n1632), .B(n1634), .CI(n1657), .CO(n1621), .S(n1622) );
  FA_X1 U1181 ( .A(n1638), .B(n1630), .CI(n1636), .CO(n1623), .S(n1624) );
  FA_X1 U1182 ( .A(n1663), .B(n1659), .CI(n1661), .CO(n1625), .S(n1626) );
  FA_X1 U1183 ( .A(n1667), .B(n1640), .CI(n1665), .CO(n1627), .S(n1628) );
  FA_X1 U1184 ( .A(n2414), .B(n2286), .CI(n2350), .CO(n1629), .S(n1630) );
  FA_X1 U1185 ( .A(n2190), .B(n2222), .CI(n2446), .CO(n1631), .S(n1632) );
  FA_X1 U1186 ( .A(n2158), .B(n2478), .CI(n2254), .CO(n1633), .S(n1634) );
  FA_X1 U1188 ( .A(n2606), .B(n2382), .CI(n2574), .CO(n1637), .S(n1638) );
  HA_X1 U1189 ( .A(n2126), .B(n2061), .CO(n1639), .S(n1640) );
  FA_X1 U1190 ( .A(n1671), .B(n1646), .CI(n1644), .CO(n1641), .S(n1642) );
  FA_X1 U1191 ( .A(n1648), .B(n1650), .CI(n1673), .CO(n1643), .S(n1644) );
  FA_X1 U1192 ( .A(n1677), .B(n1652), .CI(n1675), .CO(n1645), .S(n1646) );
  FA_X1 U1193 ( .A(n1656), .B(n1679), .CI(n1654), .CO(n1647), .S(n1648) );
  FA_X1 U1194 ( .A(n1681), .B(n1683), .CI(n1658), .CO(n1649), .S(n1650) );
  FA_X1 U1195 ( .A(n1664), .B(n1662), .CI(n1685), .CO(n1651), .S(n1652) );
  FA_X1 U1196 ( .A(n1668), .B(n1660), .CI(n1666), .CO(n1653), .S(n1654) );
  FA_X1 U1197 ( .A(n1691), .B(n1687), .CI(n1689), .CO(n1655), .S(n1656) );
  FA_X1 U1198 ( .A(n1695), .B(n2447), .CI(n1693), .CO(n1657), .S(n1658) );
  FA_X1 U1199 ( .A(n2415), .B(n2479), .CI(n2383), .CO(n1659), .S(n1660) );
  FA_X1 U1200 ( .A(n2319), .B(n2287), .CI(n2351), .CO(n1661), .S(n1662) );
  FA_X1 U1201 ( .A(n2223), .B(n2511), .CI(n2255), .CO(n1663), .S(n1664) );
  FA_X1 U1202 ( .A(n2191), .B(n2575), .CI(n2543), .CO(n1665), .S(n1666) );
  FA_X1 U1203 ( .A(n2159), .B(n2607), .CI(n2127), .CO(n1667), .S(n1668) );
  FA_X1 U1204 ( .A(n1699), .B(n1674), .CI(n1672), .CO(n1669), .S(n1670) );
  FA_X1 U1205 ( .A(n1676), .B(n1678), .CI(n1701), .CO(n1671), .S(n1672) );
  FA_X1 U1206 ( .A(n1705), .B(n1680), .CI(n1703), .CO(n1673), .S(n1674) );
  FA_X1 U1208 ( .A(n1686), .B(n1711), .CI(n1709), .CO(n1677), .S(n1678) );
  FA_X1 U1209 ( .A(n1690), .B(n1692), .CI(n1694), .CO(n1679), .S(n1680) );
  FA_X1 U1210 ( .A(n1713), .B(n1717), .CI(n1688), .CO(n1681), .S(n1682) );
  FA_X1 U1212 ( .A(n2480), .B(n2448), .CI(n1696), .CO(n1685), .S(n1686) );
  FA_X1 U1213 ( .A(n2288), .B(n2512), .CI(n2320), .CO(n1687), .S(n1688) );
  FA_X1 U1214 ( .A(n2544), .B(n2416), .CI(n2256), .CO(n1689), .S(n1690) );
  FA_X1 U1215 ( .A(n2576), .B(n2352), .CI(n2224), .CO(n1691), .S(n1692) );
  FA_X1 U1216 ( .A(n2608), .B(n2384), .CI(n2192), .CO(n1693), .S(n1694) );
  HA_X1 U1217 ( .A(n2160), .B(n2062), .CO(n1695), .S(n1696) );
  FA_X1 U1218 ( .A(n1725), .B(n1702), .CI(n1700), .CO(n1697), .S(n1698) );
  FA_X1 U1219 ( .A(n1704), .B(n1729), .CI(n1727), .CO(n1699), .S(n1700) );
  FA_X1 U1220 ( .A(n1731), .B(n1708), .CI(n1706), .CO(n1701), .S(n1702) );
  FA_X1 U1221 ( .A(n1733), .B(n1712), .CI(n1710), .CO(n1703), .S(n1704) );
  FA_X1 U1222 ( .A(n1737), .B(n1718), .CI(n1735), .CO(n1705), .S(n1706) );
  FA_X1 U1225 ( .A(n1745), .B(n1747), .CI(n1743), .CO(n1711), .S(n1712) );
  FA_X1 U1227 ( .A(n2321), .B(n2481), .CI(n2353), .CO(n1715), .S(n1716) );
  FA_X1 U1228 ( .A(n2257), .B(n2513), .CI(n2289), .CO(n1717), .S(n1718) );
  FA_X1 U1230 ( .A(n2193), .B(n2609), .CI(n2161), .CO(n1721), .S(n1722) );
  FA_X1 U1232 ( .A(n1730), .B(n1732), .CI(n1753), .CO(n1725), .S(n1726) );
  FA_X1 U1233 ( .A(n1734), .B(n1757), .CI(n1755), .CO(n1727), .S(n1728) );
  FA_X1 U1234 ( .A(n1759), .B(n1738), .CI(n1736), .CO(n1729), .S(n1730) );
  FA_X1 U1235 ( .A(n1744), .B(n1746), .CI(n1761), .CO(n1731), .S(n1732) );
  FA_X1 U1236 ( .A(n1740), .B(n1763), .CI(n1742), .CO(n1733), .S(n1734) );
  FA_X1 U1237 ( .A(n1767), .B(n1765), .CI(n1769), .CO(n1735), .S(n1736) );
  FA_X1 U1238 ( .A(n1748), .B(n2514), .CI(n1771), .CO(n1737), .S(n1738) );
  FA_X1 U1239 ( .A(n2450), .B(n2482), .CI(n2546), .CO(n1739), .S(n1740) );
  FA_X1 U1240 ( .A(n2578), .B(n2354), .CI(n2322), .CO(n1741), .S(n1742) );
  FA_X1 U1241 ( .A(n2258), .B(n2386), .CI(n2290), .CO(n1743), .S(n1744) );
  FA_X1 U1242 ( .A(n2226), .B(n2418), .CI(n2610), .CO(n1745), .S(n1746) );
  HA_X1 U1243 ( .A(n2194), .B(n2063), .CO(n1747), .S(n1748) );
  FA_X1 U1244 ( .A(n1775), .B(n1754), .CI(n1752), .CO(n1749), .S(n1750) );
  FA_X1 U1245 ( .A(n1777), .B(n1779), .CI(n1756), .CO(n1751), .S(n1752) );
  FA_X1 U1246 ( .A(n1760), .B(n1762), .CI(n1758), .CO(n1753), .S(n1754) );
  FA_X1 U1247 ( .A(n1783), .B(n1785), .CI(n1781), .CO(n1755), .S(n1756) );
  FA_X1 U1248 ( .A(n1770), .B(n1772), .CI(n1764), .CO(n1757), .S(n1758) );
  FA_X1 U1249 ( .A(n1766), .B(n1793), .CI(n1768), .CO(n1759), .S(n1760) );
  FA_X1 U1250 ( .A(n1787), .B(n1789), .CI(n1791), .CO(n1761), .S(n1762) );
  FA_X1 U1251 ( .A(n2451), .B(n2483), .CI(n1795), .CO(n1763), .S(n1764) );
  FA_X1 U1252 ( .A(n2387), .B(n2515), .CI(n2419), .CO(n1765), .S(n1766) );
  FA_X1 U1254 ( .A(n2259), .B(n2579), .CI(n2291), .CO(n1769), .S(n1770) );
  FA_X1 U1255 ( .A(n2227), .B(n2611), .CI(n2195), .CO(n1771), .S(n1772) );
  FA_X1 U1257 ( .A(n1780), .B(n1803), .CI(n1801), .CO(n1775), .S(n1776) );
  FA_X1 U1258 ( .A(n1784), .B(n1805), .CI(n1782), .CO(n1777), .S(n1778) );
  FA_X1 U1259 ( .A(n1807), .B(n1809), .CI(n1786), .CO(n1779), .S(n1780) );
  FA_X1 U1260 ( .A(n1794), .B(n1790), .CI(n1792), .CO(n1781), .S(n1782) );
  FA_X1 U1261 ( .A(n1811), .B(n1813), .CI(n1788), .CO(n1783), .S(n1784) );
  FA_X1 U1262 ( .A(n1817), .B(n1796), .CI(n1815), .CO(n1785), .S(n1786) );
  FA_X1 U1263 ( .A(n2356), .B(n2484), .CI(n2452), .CO(n1787), .S(n1788) );
  FA_X1 U1264 ( .A(n2292), .B(n2516), .CI(n2324), .CO(n1789), .S(n1790) );
  FA_X1 U1265 ( .A(n2580), .B(n2388), .CI(n2548), .CO(n1791), .S(n1792) );
  FA_X1 U1266 ( .A(n2612), .B(n2420), .CI(n2260), .CO(n1793), .S(n1794) );
  HA_X1 U1267 ( .A(n2228), .B(n2064), .CO(n1795), .S(n1796) );
  FA_X1 U1269 ( .A(n1804), .B(n1825), .CI(n1823), .CO(n1799), .S(n1800) );
  FA_X1 U1270 ( .A(n1808), .B(n1827), .CI(n1806), .CO(n1801), .S(n1802) );
  FA_X1 U1271 ( .A(n1829), .B(n1831), .CI(n1810), .CO(n1803), .S(n1804) );
  FA_X1 U1272 ( .A(n1818), .B(n1814), .CI(n1816), .CO(n1805), .S(n1806) );
  FA_X1 U1273 ( .A(n1833), .B(n1835), .CI(n1812), .CO(n1807), .S(n1808) );
  FA_X1 U1274 ( .A(n1839), .B(n2453), .CI(n1837), .CO(n1809), .S(n1810) );
  FA_X1 U1275 ( .A(n2389), .B(n2421), .CI(n2485), .CO(n1811), .S(n1812) );
  FA_X1 U1276 ( .A(n2357), .B(n2549), .CI(n2517), .CO(n1813), .S(n1814) );
  FA_X1 U1277 ( .A(n2293), .B(n2581), .CI(n2325), .CO(n1815), .S(n1816) );
  FA_X1 U1278 ( .A(n2261), .B(n2613), .CI(n2229), .CO(n1817), .S(n1818) );
  FA_X1 U1279 ( .A(n1843), .B(n1824), .CI(n1822), .CO(n1819), .S(n1820) );
  FA_X1 U1280 ( .A(n1845), .B(n1828), .CI(n1826), .CO(n1821), .S(n1822) );
  FA_X1 U1281 ( .A(n1830), .B(n1849), .CI(n1847), .CO(n1823), .S(n1824) );
  FA_X1 U1282 ( .A(n1851), .B(n1838), .CI(n1832), .CO(n1825), .S(n1826) );
  FA_X1 U1283 ( .A(n1834), .B(n1857), .CI(n1836), .CO(n1827), .S(n1828) );
  FA_X1 U1284 ( .A(n1853), .B(n1859), .CI(n1855), .CO(n1829), .S(n1830) );
  FA_X1 U1285 ( .A(n2486), .B(n2518), .CI(n1840), .CO(n1831), .S(n1832) );
  FA_X1 U1286 ( .A(n2358), .B(n2550), .CI(n2390), .CO(n1833), .S(n1834) );
  FA_X1 U1287 ( .A(n2582), .B(n2422), .CI(n2326), .CO(n1835), .S(n1836) );
  FA_X1 U1288 ( .A(n2614), .B(n2454), .CI(n2294), .CO(n1837), .S(n1838) );
  HA_X1 U1289 ( .A(n2262), .B(n2065), .CO(n1839), .S(n1840) );
  FA_X1 U1290 ( .A(n1863), .B(n1846), .CI(n1844), .CO(n1841), .S(n1842) );
  FA_X1 U1291 ( .A(n1848), .B(n1850), .CI(n1865), .CO(n1843), .S(n1844) );
  FA_X1 U1292 ( .A(n1852), .B(n1869), .CI(n1867), .CO(n1845), .S(n1846) );
  FA_X1 U1293 ( .A(n1860), .B(n1858), .CI(n1871), .CO(n1847), .S(n1848) );
  FA_X1 U1294 ( .A(n1854), .B(n1873), .CI(n1856), .CO(n1849), .S(n1850) );
  FA_X1 U1295 ( .A(n1877), .B(n1879), .CI(n1875), .CO(n1851), .S(n1852) );
  FA_X1 U1296 ( .A(n2455), .B(n2519), .CI(n2487), .CO(n1853), .S(n1854) );
  FA_X1 U1297 ( .A(n2391), .B(n2551), .CI(n2423), .CO(n1855), .S(n1856) );
  FA_X1 U1298 ( .A(n2327), .B(n2583), .CI(n2359), .CO(n1857), .S(n1858) );
  FA_X1 U1299 ( .A(n2295), .B(n2615), .CI(n2263), .CO(n1859), .S(n1860) );
  FA_X1 U1300 ( .A(n1883), .B(n1866), .CI(n1864), .CO(n1861), .S(n1862) );
  FA_X1 U1301 ( .A(n1868), .B(n1870), .CI(n1885), .CO(n1863), .S(n1864) );
  FA_X1 U1302 ( .A(n1872), .B(n1889), .CI(n1887), .CO(n1865), .S(n1866) );
  FA_X1 U1303 ( .A(n1878), .B(n1874), .CI(n1876), .CO(n1867), .S(n1868) );
  FA_X1 U1304 ( .A(n1893), .B(n1895), .CI(n1891), .CO(n1869), .S(n1870) );
  FA_X1 U1305 ( .A(n1880), .B(n2488), .CI(n1897), .CO(n1871), .S(n1872) );
  FA_X1 U1306 ( .A(n2360), .B(n2520), .CI(n2392), .CO(n1873), .S(n1874) );
  FA_X1 U1307 ( .A(n2328), .B(n2424), .CI(n2552), .CO(n1875), .S(n1876) );
  FA_X1 U1308 ( .A(n2616), .B(n2584), .CI(n2456), .CO(n1877), .S(n1878) );
  HA_X1 U1309 ( .A(n2296), .B(n2066), .CO(n1879), .S(n1880) );
  FA_X1 U1310 ( .A(n1901), .B(n1886), .CI(n1884), .CO(n1881), .S(n1882) );
  FA_X1 U1311 ( .A(n1888), .B(n1890), .CI(n1903), .CO(n1883), .S(n1884) );
  FA_X1 U1312 ( .A(n1907), .B(n1892), .CI(n1905), .CO(n1885), .S(n1886) );
  FA_X1 U1313 ( .A(n1898), .B(n1894), .CI(n1896), .CO(n1887), .S(n1888) );
  FA_X1 U1314 ( .A(n1909), .B(n1913), .CI(n1911), .CO(n1889), .S(n1890) );
  FA_X1 U1315 ( .A(n2489), .B(n2521), .CI(n1915), .CO(n1891), .S(n1892) );
  FA_X1 U1316 ( .A(n2425), .B(n2553), .CI(n2457), .CO(n1893), .S(n1894) );
  FA_X1 U1317 ( .A(n2361), .B(n2585), .CI(n2393), .CO(n1895), .S(n1896) );
  FA_X1 U1318 ( .A(n2297), .B(n2617), .CI(n2329), .CO(n1897), .S(n1898) );
  FA_X1 U1319 ( .A(n1919), .B(n1904), .CI(n1902), .CO(n1899), .S(n1900) );
  FA_X1 U1320 ( .A(n1906), .B(n1923), .CI(n1921), .CO(n1901), .S(n1902) );
  FA_X1 U1321 ( .A(n1925), .B(n1914), .CI(n1908), .CO(n1903), .S(n1904) );
  FA_X1 U1322 ( .A(n1910), .B(n1927), .CI(n1912), .CO(n1905), .S(n1906) );
  FA_X1 U1323 ( .A(n1931), .B(n1916), .CI(n1929), .CO(n1907), .S(n1908) );
  FA_X1 U1324 ( .A(n2458), .B(n2586), .CI(n2554), .CO(n1909), .S(n1910) );
  FA_X1 U1325 ( .A(n2618), .B(n2522), .CI(n2426), .CO(n1911), .S(n1912) );
  FA_X1 U1326 ( .A(n2362), .B(n2490), .CI(n2394), .CO(n1913), .S(n1914) );
  HA_X1 U1327 ( .A(n2330), .B(n2067), .CO(n1915), .S(n1916) );
  FA_X1 U1328 ( .A(n1935), .B(n1922), .CI(n1920), .CO(n1917), .S(n1918) );
  FA_X1 U1329 ( .A(n1924), .B(n1926), .CI(n1937), .CO(n1919), .S(n1920) );
  FA_X1 U1330 ( .A(n1941), .B(n1932), .CI(n1939), .CO(n1921), .S(n1922) );
  FA_X1 U1331 ( .A(n1928), .B(n1943), .CI(n1930), .CO(n1923), .S(n1924) );
  FA_X1 U1332 ( .A(n1947), .B(n2523), .CI(n1945), .CO(n1925), .S(n1926) );
  FA_X1 U1333 ( .A(n2459), .B(n2491), .CI(n2555), .CO(n1927), .S(n1928) );
  FA_X1 U1334 ( .A(n2427), .B(n2587), .CI(n2395), .CO(n1929), .S(n1930) );
  FA_X1 U1335 ( .A(n2363), .B(n2619), .CI(n2331), .CO(n1931), .S(n1932) );
  FA_X1 U1336 ( .A(n1938), .B(n1951), .CI(n1936), .CO(n1933), .S(n1934) );
  FA_X1 U1337 ( .A(n1953), .B(n1942), .CI(n1940), .CO(n1935), .S(n1936) );
  FA_X1 U1338 ( .A(n1946), .B(n1944), .CI(n1955), .CO(n1937), .S(n1938) );
  FA_X1 U1339 ( .A(n1957), .B(n1961), .CI(n1959), .CO(n1939), .S(n1940) );
  FA_X1 U1340 ( .A(n2556), .B(n2588), .CI(n1948), .CO(n1941), .S(n1942) );
  FA_X1 U1341 ( .A(n2428), .B(n2524), .CI(n2460), .CO(n1943), .S(n1944) );
  FA_X1 U1342 ( .A(n2396), .B(n2492), .CI(n2620), .CO(n1945), .S(n1946) );
  HA_X1 U1343 ( .A(n2364), .B(n2068), .CO(n1947), .S(n1948) );
  FA_X1 U1344 ( .A(n1965), .B(n1954), .CI(n1952), .CO(n1949), .S(n1950) );
  FA_X1 U1345 ( .A(n1967), .B(n1969), .CI(n1956), .CO(n1951), .S(n1952) );
  FA_X1 U1346 ( .A(n1960), .B(n1962), .CI(n1958), .CO(n1953), .S(n1954) );
  FA_X1 U1347 ( .A(n1973), .B(n1975), .CI(n1971), .CO(n1955), .S(n1956) );
  FA_X1 U1348 ( .A(n2493), .B(n2557), .CI(n2525), .CO(n1957), .S(n1958) );
  FA_X1 U1349 ( .A(n2429), .B(n2589), .CI(n2461), .CO(n1959), .S(n1960) );
  FA_X1 U1350 ( .A(n2397), .B(n2621), .CI(n2365), .CO(n1961), .S(n1962) );
  FA_X1 U1351 ( .A(n1979), .B(n1968), .CI(n1966), .CO(n1963), .S(n1964) );
  FA_X1 U1352 ( .A(n1981), .B(n1974), .CI(n1970), .CO(n1965), .S(n1966) );
  FA_X1 U1353 ( .A(n1983), .B(n1985), .CI(n1972), .CO(n1967), .S(n1968) );
  FA_X1 U1354 ( .A(n1976), .B(n2494), .CI(n1987), .CO(n1969), .S(n1970) );
  FA_X1 U1355 ( .A(n2558), .B(n2430), .CI(n2462), .CO(n1971), .S(n1972) );
  FA_X1 U1356 ( .A(n2622), .B(n2526), .CI(n2590), .CO(n1973), .S(n1974) );
  HA_X1 U1357 ( .A(n2398), .B(n2069), .CO(n1975), .S(n1976) );
  FA_X1 U1358 ( .A(n1991), .B(n1982), .CI(n1980), .CO(n1977), .S(n1978) );
  FA_X1 U1359 ( .A(n1984), .B(n1988), .CI(n1993), .CO(n1979), .S(n1980) );
  FA_X1 U1360 ( .A(n1995), .B(n1997), .CI(n1986), .CO(n1981), .S(n1982) );
  FA_X1 U1361 ( .A(n2527), .B(n2559), .CI(n1999), .CO(n1983), .S(n1984) );
  FA_X1 U1362 ( .A(n2463), .B(n2591), .CI(n2495), .CO(n1985), .S(n1986) );
  FA_X1 U1363 ( .A(n2431), .B(n2623), .CI(n2399), .CO(n1987), .S(n1988) );
  FA_X1 U1364 ( .A(n2003), .B(n1994), .CI(n1992), .CO(n1989), .S(n1990) );
  FA_X1 U1365 ( .A(n1998), .B(n1996), .CI(n2005), .CO(n1991), .S(n1992) );
  FA_X1 U1366 ( .A(n2009), .B(n2000), .CI(n2007), .CO(n1993), .S(n1994) );
  FA_X1 U1367 ( .A(n2464), .B(n2560), .CI(n2496), .CO(n1995), .S(n1996) );
  FA_X1 U1368 ( .A(n2624), .B(n2528), .CI(n2592), .CO(n1997), .S(n1998) );
  HA_X1 U1369 ( .A(n2432), .B(n2070), .CO(n1999), .S(n2000) );
  FA_X1 U1370 ( .A(n2006), .B(n2013), .CI(n2004), .CO(n2001), .S(n2002) );
  FA_X1 U1371 ( .A(n2010), .B(n2008), .CI(n2015), .CO(n2003), .S(n2004) );
  FA_X1 U1372 ( .A(n2019), .B(n2561), .CI(n2017), .CO(n2005), .S(n2006) );
  FA_X1 U1373 ( .A(n2497), .B(n2593), .CI(n2529), .CO(n2007), .S(n2008) );
  FA_X1 U1374 ( .A(n2465), .B(n2625), .CI(n2433), .CO(n2009), .S(n2010) );
  FA_X1 U1375 ( .A(n2023), .B(n2016), .CI(n2014), .CO(n2011), .S(n2012) );
  FA_X1 U1376 ( .A(n2025), .B(n2027), .CI(n2018), .CO(n2013), .S(n2014) );
  FA_X1 U1377 ( .A(n2498), .B(n2530), .CI(n2020), .CO(n2015), .S(n2016) );
  FA_X1 U1378 ( .A(n2626), .B(n2562), .CI(n2594), .CO(n2017), .S(n2018) );
  HA_X1 U1379 ( .A(n2466), .B(n2071), .CO(n2019), .S(n2020) );
  FA_X1 U1380 ( .A(n2031), .B(n2028), .CI(n2024), .CO(n2021), .S(n2022) );
  FA_X1 U1381 ( .A(n2033), .B(n2035), .CI(n2026), .CO(n2023), .S(n2024) );
  FA_X1 U1382 ( .A(n2531), .B(n2595), .CI(n2563), .CO(n2025), .S(n2026) );
  FA_X1 U1383 ( .A(n2499), .B(n2627), .CI(n2467), .CO(n2027), .S(n2028) );
  FA_X1 U1384 ( .A(n2034), .B(n2039), .CI(n2032), .CO(n2029), .S(n2030) );
  FA_X1 U1385 ( .A(n2036), .B(n2628), .CI(n2041), .CO(n2031), .S(n2032) );
  FA_X1 U1386 ( .A(n2532), .B(n2564), .CI(n2596), .CO(n2033), .S(n2034) );
  HA_X1 U1387 ( .A(n2500), .B(n2072), .CO(n2035), .S(n2036) );
  FA_X1 U1388 ( .A(n2042), .B(n2045), .CI(n2040), .CO(n2037), .S(n2038) );
  FA_X1 U1389 ( .A(n2565), .B(n2597), .CI(n2047), .CO(n2039), .S(n2040) );
  FA_X1 U1390 ( .A(n2533), .B(n2629), .CI(n2501), .CO(n2041), .S(n2042) );
  FA_X1 U1391 ( .A(n2051), .B(n2048), .CI(n2046), .CO(n2043), .S(n2044) );
  FA_X1 U1392 ( .A(n2566), .B(n2630), .CI(n2598), .CO(n2045), .S(n2046) );
  HA_X1 U1393 ( .A(n2534), .B(n2073), .CO(n2047), .S(n2048) );
  FA_X1 U1394 ( .A(n2055), .B(n2599), .CI(n2052), .CO(n2049), .S(n2050) );
  FA_X1 U1395 ( .A(n2567), .B(n2631), .CI(n2535), .CO(n2051), .S(n2052) );
  FA_X1 U1396 ( .A(n2600), .B(n2632), .CI(n2056), .CO(n2053), .S(n2054) );
  HA_X1 U1397 ( .A(n2568), .B(n2074), .CO(n2055), .S(n2056) );
  FA_X1 U1398 ( .A(n2601), .B(n2633), .CI(n2569), .CO(n2057), .S(n2058) );
  HA_X1 U1399 ( .A(n2634), .B(n2602), .CO(n2059), .S(n2060) );
  NOR2_X4 U1400 ( .A1(n2637), .A2(n3500), .ZN(n2077) );
  NOR2_X4 U1401 ( .A1(n2638), .A2(n3500), .ZN(n1044) );
  NOR2_X4 U1402 ( .A1(n2639), .A2(n3500), .ZN(n2078) );
  NOR2_X4 U1403 ( .A1(n2640), .A2(n3500), .ZN(n1054) );
  NOR2_X4 U1404 ( .A1(n2641), .A2(n3500), .ZN(n2079) );
  NOR2_X4 U1405 ( .A1(n2642), .A2(n3500), .ZN(n1068) );
  NOR2_X4 U1406 ( .A1(n2643), .A2(n3500), .ZN(n2080) );
  NOR2_X4 U1407 ( .A1(n2644), .A2(n3500), .ZN(n1086) );
  NOR2_X4 U1408 ( .A1(n2645), .A2(n3500), .ZN(n2081) );
  NOR2_X4 U1409 ( .A1(n2646), .A2(n3500), .ZN(n1108) );
  NOR2_X4 U1410 ( .A1(n2647), .A2(n3500), .ZN(n2082) );
  NOR2_X4 U1411 ( .A1(n2648), .A2(n3500), .ZN(n1134) );
  NOR2_X4 U1412 ( .A1(n2649), .A2(n3500), .ZN(n2083) );
  NOR2_X4 U1413 ( .A1(n2650), .A2(n3500), .ZN(n1164) );
  NOR2_X4 U1414 ( .A1(n2651), .A2(n3500), .ZN(n2084) );
  NOR2_X4 U1415 ( .A1(n2652), .A2(n3500), .ZN(n1198) );
  NOR2_X4 U1416 ( .A1(n2653), .A2(n3500), .ZN(n2085) );
  NOR2_X4 U1417 ( .A1(n2654), .A2(n3500), .ZN(n1236) );
  NOR2_X4 U1418 ( .A1(n2655), .A2(n3500), .ZN(n2086) );
  NOR2_X4 U1419 ( .A1(n2656), .A2(n3500), .ZN(n1278) );
  NOR2_X4 U1420 ( .A1(n2657), .A2(n3500), .ZN(n2087) );
  NOR2_X4 U1421 ( .A1(n2658), .A2(n3500), .ZN(n1324) );
  NOR2_X4 U1422 ( .A1(n2659), .A2(n3500), .ZN(n2088) );
  NOR2_X4 U1423 ( .A1(n2660), .A2(n3500), .ZN(n1374) );
  NOR2_X4 U1424 ( .A1(n2661), .A2(n3500), .ZN(n2089) );
  NOR2_X4 U1425 ( .A1(n2662), .A2(n3500), .ZN(n1428) );
  NOR2_X4 U1426 ( .A1(n2663), .A2(n3500), .ZN(n2090) );
  NOR2_X4 U1427 ( .A1(n2664), .A2(n3500), .ZN(n1486) );
  NOR2_X4 U1428 ( .A1(n2665), .A2(n3500), .ZN(n2091) );
  NOR2_X4 U1429 ( .A1(n2666), .A2(n3500), .ZN(n2092) );
  NOR2_X4 U1430 ( .A1(n2667), .A2(n3500), .ZN(n1548) );
  OAI22_X2 U1463 ( .A1(n3653), .A2(n2668), .B1(n3625), .B2(n3500), .ZN(n2095)
         );
  OAI22_X2 U1465 ( .A1(n3653), .A2(n2670), .B1(n2669), .B2(n3625), .ZN(n2097)
         );
  OAI22_X2 U1466 ( .A1(n3653), .A2(n2671), .B1(n2670), .B2(n3625), .ZN(n2098)
         );
  OAI22_X2 U1592 ( .A1(n458), .A2(n3279), .B1(n2766), .B2(n3638), .ZN(n2063)
         );
  OAI22_X2 U1593 ( .A1(n458), .A2(n2734), .B1(n3638), .B2(n3279), .ZN(n2163)
         );
  OAI22_X2 U1594 ( .A1(n458), .A2(n2735), .B1(n2734), .B2(n3639), .ZN(n2164)
         );
  OAI22_X2 U1595 ( .A1(n458), .A2(n2736), .B1(n2735), .B2(n3639), .ZN(n2165)
         );
  OAI22_X2 U1596 ( .A1(n458), .A2(n2737), .B1(n2736), .B2(n3638), .ZN(n2166)
         );
  OAI22_X2 U1597 ( .A1(n458), .A2(n2738), .B1(n2737), .B2(n3638), .ZN(n2167)
         );
  OAI22_X2 U1598 ( .A1(n458), .A2(n2739), .B1(n2738), .B2(n3639), .ZN(n2168)
         );
  OAI22_X2 U1599 ( .A1(n458), .A2(n2740), .B1(n2739), .B2(n3638), .ZN(n2169)
         );
  OAI22_X2 U1600 ( .A1(n458), .A2(n2741), .B1(n2740), .B2(n3638), .ZN(n2170)
         );
  OAI22_X2 U1601 ( .A1(n458), .A2(n2742), .B1(n2741), .B2(n3639), .ZN(n2171)
         );
  OAI22_X2 U1602 ( .A1(n458), .A2(n2743), .B1(n2742), .B2(n3638), .ZN(n2172)
         );
  OAI22_X2 U1603 ( .A1(n458), .A2(n2744), .B1(n2743), .B2(n3638), .ZN(n2173)
         );
  OAI22_X2 U1604 ( .A1(n458), .A2(n2745), .B1(n2744), .B2(n3639), .ZN(n2174)
         );
  OAI22_X2 U1605 ( .A1(n458), .A2(n2746), .B1(n2745), .B2(n3638), .ZN(n2175)
         );
  OAI22_X2 U1606 ( .A1(n458), .A2(n2747), .B1(n2746), .B2(n3639), .ZN(n2176)
         );
  OAI22_X2 U1607 ( .A1(n458), .A2(n2748), .B1(n2747), .B2(n3638), .ZN(n2177)
         );
  OAI22_X2 U1608 ( .A1(n458), .A2(n2749), .B1(n2748), .B2(n3639), .ZN(n2178)
         );
  OAI22_X2 U1609 ( .A1(n458), .A2(n2750), .B1(n2749), .B2(n3639), .ZN(n2179)
         );
  OAI22_X2 U1610 ( .A1(n458), .A2(n2751), .B1(n2750), .B2(n3638), .ZN(n2180)
         );
  OAI22_X2 U1611 ( .A1(n458), .A2(n2752), .B1(n2751), .B2(n3639), .ZN(n2181)
         );
  OAI22_X2 U1612 ( .A1(n458), .A2(n2753), .B1(n2752), .B2(n3639), .ZN(n2182)
         );
  OAI22_X2 U1613 ( .A1(n458), .A2(n2754), .B1(n2753), .B2(n3639), .ZN(n2183)
         );
  OAI22_X2 U1614 ( .A1(n458), .A2(n2755), .B1(n2754), .B2(n3638), .ZN(n2184)
         );
  OAI22_X2 U1615 ( .A1(n458), .A2(n2756), .B1(n2755), .B2(n3639), .ZN(n2185)
         );
  OAI22_X2 U1616 ( .A1(n458), .A2(n2757), .B1(n2756), .B2(n3638), .ZN(n2186)
         );
  OAI22_X2 U1619 ( .A1(n458), .A2(n2760), .B1(n2759), .B2(n3638), .ZN(n2189)
         );
  OAI22_X2 U1621 ( .A1(n458), .A2(n2762), .B1(n2761), .B2(n3639), .ZN(n2191)
         );
  OAI22_X2 U1623 ( .A1(n458), .A2(n2764), .B1(n2763), .B2(n3639), .ZN(n2193)
         );
  OAI22_X2 U1624 ( .A1(n458), .A2(n2765), .B1(n2764), .B2(n3639), .ZN(n2194)
         );
  OAI22_X2 U1659 ( .A1(n3462), .A2(n2768), .B1(n2767), .B2(n405), .ZN(n2198)
         );
  OAI22_X2 U1660 ( .A1(n3461), .A2(n2769), .B1(n2768), .B2(n405), .ZN(n2199)
         );
  OAI22_X2 U1661 ( .A1(n3462), .A2(n2770), .B1(n2769), .B2(n405), .ZN(n2200)
         );
  OAI22_X2 U1662 ( .A1(n3461), .A2(n2771), .B1(n2770), .B2(n405), .ZN(n2201)
         );
  OAI22_X2 U1663 ( .A1(n3461), .A2(n2772), .B1(n2771), .B2(n405), .ZN(n2202)
         );
  OAI22_X2 U1664 ( .A1(n3462), .A2(n2773), .B1(n2772), .B2(n405), .ZN(n2203)
         );
  OAI22_X2 U1665 ( .A1(n3461), .A2(n2774), .B1(n2773), .B2(n405), .ZN(n2204)
         );
  OAI22_X2 U1666 ( .A1(n3462), .A2(n2775), .B1(n2774), .B2(n405), .ZN(n2205)
         );
  OAI22_X2 U1667 ( .A1(n3462), .A2(n2776), .B1(n2775), .B2(n405), .ZN(n2206)
         );
  OAI22_X2 U1668 ( .A1(n3461), .A2(n2777), .B1(n2776), .B2(n405), .ZN(n2207)
         );
  OAI22_X2 U1669 ( .A1(n3462), .A2(n2778), .B1(n2777), .B2(n405), .ZN(n2208)
         );
  OAI22_X2 U1670 ( .A1(n3462), .A2(n2779), .B1(n2778), .B2(n405), .ZN(n2209)
         );
  OAI22_X2 U1671 ( .A1(n3461), .A2(n2780), .B1(n2779), .B2(n405), .ZN(n2210)
         );
  OAI22_X2 U1672 ( .A1(n3461), .A2(n2781), .B1(n2780), .B2(n405), .ZN(n2211)
         );
  OAI22_X2 U1673 ( .A1(n3461), .A2(n2782), .B1(n2781), .B2(n405), .ZN(n2212)
         );
  OAI22_X2 U1674 ( .A1(n3462), .A2(n2783), .B1(n2782), .B2(n405), .ZN(n2213)
         );
  OAI22_X2 U1675 ( .A1(n3461), .A2(n2784), .B1(n2783), .B2(n405), .ZN(n2214)
         );
  OAI22_X2 U1676 ( .A1(n3462), .A2(n2785), .B1(n2784), .B2(n405), .ZN(n2215)
         );
  OAI22_X2 U1677 ( .A1(n3461), .A2(n2786), .B1(n2785), .B2(n405), .ZN(n2216)
         );
  OAI22_X2 U1678 ( .A1(n3461), .A2(n2787), .B1(n2786), .B2(n405), .ZN(n2217)
         );
  OAI22_X2 U1681 ( .A1(n3462), .A2(n2790), .B1(n2789), .B2(n405), .ZN(n2220)
         );
  OAI22_X2 U1682 ( .A1(n3461), .A2(n2791), .B1(n2790), .B2(n405), .ZN(n2221)
         );
  OAI22_X2 U1683 ( .A1(n3462), .A2(n2792), .B1(n2791), .B2(n405), .ZN(n2222)
         );
  OAI22_X2 U1684 ( .A1(n3461), .A2(n2793), .B1(n2792), .B2(n405), .ZN(n2223)
         );
  OAI22_X2 U1685 ( .A1(n3462), .A2(n2794), .B1(n2793), .B2(n405), .ZN(n2224)
         );
  OAI22_X2 U1687 ( .A1(n3462), .A2(n2796), .B1(n2795), .B2(n405), .ZN(n2226)
         );
  OAI22_X2 U1688 ( .A1(n3462), .A2(n2797), .B1(n2796), .B2(n405), .ZN(n2227)
         );
  OAI22_X2 U1689 ( .A1(n3462), .A2(n2798), .B1(n2797), .B2(n405), .ZN(n2228)
         );
  OAI22_X2 U1787 ( .A1(n3643), .A2(n3282), .B1(n2865), .B2(n399), .ZN(n2066)
         );
  OAI22_X2 U1788 ( .A1(n3643), .A2(n2833), .B1(n399), .B2(n3282), .ZN(n2265)
         );
  OAI22_X2 U1790 ( .A1(n3643), .A2(n2835), .B1(n2834), .B2(n399), .ZN(n2267)
         );
  OAI22_X2 U1793 ( .A1(n3643), .A2(n2838), .B1(n2837), .B2(n399), .ZN(n2270)
         );
  OAI22_X2 U1794 ( .A1(n3643), .A2(n2839), .B1(n2838), .B2(n399), .ZN(n2271)
         );
  OAI22_X2 U1797 ( .A1(n3643), .A2(n2842), .B1(n2841), .B2(n399), .ZN(n2274)
         );
  OAI22_X2 U1798 ( .A1(n3643), .A2(n2843), .B1(n2842), .B2(n399), .ZN(n2275)
         );
  OAI22_X2 U1802 ( .A1(n3643), .A2(n2847), .B1(n2846), .B2(n399), .ZN(n2279)
         );
  OAI22_X2 U1807 ( .A1(n3643), .A2(n2852), .B1(n2851), .B2(n399), .ZN(n2284)
         );
  OAI22_X2 U1811 ( .A1(n3643), .A2(n2856), .B1(n2855), .B2(n399), .ZN(n2288)
         );
  OAI22_X2 U1813 ( .A1(n3643), .A2(n2858), .B1(n2857), .B2(n399), .ZN(n2290)
         );
  OAI22_X2 U1814 ( .A1(n3643), .A2(n2859), .B1(n2858), .B2(n399), .ZN(n2291)
         );
  OAI22_X2 U1816 ( .A1(n3643), .A2(n2861), .B1(n2860), .B2(n399), .ZN(n2293)
         );
  OAI22_X2 U1818 ( .A1(n3643), .A2(n2863), .B1(n2862), .B2(n399), .ZN(n2295)
         );
  OAI22_X2 U1819 ( .A1(n3643), .A2(n2864), .B1(n2863), .B2(n399), .ZN(n2296)
         );
  OAI22_X2 U1917 ( .A1(n443), .A2(n3284), .B1(n2931), .B2(n3656), .ZN(n2068)
         );
  OAI22_X2 U1918 ( .A1(n443), .A2(n2899), .B1(n3656), .B2(n3284), .ZN(n2333)
         );
  OAI22_X2 U1919 ( .A1(n443), .A2(n2900), .B1(n2899), .B2(n3656), .ZN(n2334)
         );
  OAI22_X2 U1920 ( .A1(n443), .A2(n2901), .B1(n2900), .B2(n3656), .ZN(n2335)
         );
  OAI22_X2 U1921 ( .A1(n443), .A2(n2902), .B1(n2901), .B2(n3656), .ZN(n2336)
         );
  OAI22_X2 U1922 ( .A1(n443), .A2(n2903), .B1(n2902), .B2(n3656), .ZN(n2337)
         );
  OAI22_X2 U1923 ( .A1(n443), .A2(n2904), .B1(n2903), .B2(n3656), .ZN(n2338)
         );
  OAI22_X2 U1924 ( .A1(n443), .A2(n2905), .B1(n2904), .B2(n3656), .ZN(n2339)
         );
  OAI22_X2 U1925 ( .A1(n443), .A2(n2906), .B1(n2905), .B2(n3656), .ZN(n2340)
         );
  OAI22_X2 U1926 ( .A1(n443), .A2(n2907), .B1(n2906), .B2(n3656), .ZN(n2341)
         );
  OAI22_X2 U1927 ( .A1(n443), .A2(n2908), .B1(n2907), .B2(n3656), .ZN(n2342)
         );
  OAI22_X2 U1928 ( .A1(n443), .A2(n2909), .B1(n2908), .B2(n3656), .ZN(n2343)
         );
  OAI22_X2 U1929 ( .A1(n443), .A2(n2910), .B1(n2909), .B2(n3656), .ZN(n2344)
         );
  OAI22_X2 U1930 ( .A1(n443), .A2(n2911), .B1(n2910), .B2(n3656), .ZN(n2345)
         );
  OAI22_X2 U1931 ( .A1(n443), .A2(n2912), .B1(n2911), .B2(n3656), .ZN(n2346)
         );
  OAI22_X2 U1932 ( .A1(n443), .A2(n2913), .B1(n2912), .B2(n3656), .ZN(n2347)
         );
  OAI22_X2 U1934 ( .A1(n443), .A2(n2915), .B1(n2914), .B2(n3656), .ZN(n2349)
         );
  OAI22_X2 U1935 ( .A1(n443), .A2(n2916), .B1(n2915), .B2(n3656), .ZN(n2350)
         );
  OAI22_X2 U1936 ( .A1(n443), .A2(n2917), .B1(n2916), .B2(n3656), .ZN(n2351)
         );
  OAI22_X2 U1937 ( .A1(n443), .A2(n2918), .B1(n2917), .B2(n3656), .ZN(n2352)
         );
  OAI22_X2 U1938 ( .A1(n443), .A2(n2919), .B1(n2918), .B2(n3656), .ZN(n2353)
         );
  OAI22_X2 U1939 ( .A1(n443), .A2(n2920), .B1(n2919), .B2(n3656), .ZN(n2354)
         );
  OAI22_X2 U1941 ( .A1(n443), .A2(n2922), .B1(n2921), .B2(n3656), .ZN(n2356)
         );
  OAI22_X2 U1942 ( .A1(n443), .A2(n2923), .B1(n2922), .B2(n3656), .ZN(n2357)
         );
  OAI22_X2 U1943 ( .A1(n443), .A2(n2924), .B1(n2923), .B2(n3656), .ZN(n2358)
         );
  OAI22_X2 U1944 ( .A1(n443), .A2(n2925), .B1(n2924), .B2(n3656), .ZN(n2359)
         );
  OAI22_X2 U1945 ( .A1(n443), .A2(n2926), .B1(n2925), .B2(n3656), .ZN(n2360)
         );
  OAI22_X2 U1946 ( .A1(n443), .A2(n2927), .B1(n2926), .B2(n3656), .ZN(n2361)
         );
  OAI22_X2 U1947 ( .A1(n443), .A2(n2928), .B1(n2927), .B2(n3656), .ZN(n2362)
         );
  OAI22_X2 U1948 ( .A1(n443), .A2(n2929), .B1(n2928), .B2(n3656), .ZN(n2363)
         );
  OAI22_X2 U1949 ( .A1(n443), .A2(n2930), .B1(n2929), .B2(n3656), .ZN(n2364)
         );
  OAI22_X2 U2047 ( .A1(n3416), .A2(n3286), .B1(n2997), .B2(n387), .ZN(n2070)
         );
  OAI22_X2 U2048 ( .A1(n3416), .A2(n2965), .B1(n387), .B2(n3286), .ZN(n2401)
         );
  OAI22_X2 U2049 ( .A1(n3416), .A2(n2966), .B1(n2965), .B2(n387), .ZN(n2402)
         );
  OAI22_X2 U2050 ( .A1(n3416), .A2(n2967), .B1(n2966), .B2(n387), .ZN(n2403)
         );
  OAI22_X2 U2051 ( .A1(n3416), .A2(n2968), .B1(n2967), .B2(n387), .ZN(n2404)
         );
  OAI22_X2 U2052 ( .A1(n3416), .A2(n2969), .B1(n2968), .B2(n387), .ZN(n2405)
         );
  OAI22_X2 U2053 ( .A1(n3416), .A2(n2970), .B1(n2969), .B2(n387), .ZN(n2406)
         );
  OAI22_X2 U2054 ( .A1(n3416), .A2(n2971), .B1(n2970), .B2(n387), .ZN(n2407)
         );
  OAI22_X2 U2055 ( .A1(n3416), .A2(n2972), .B1(n2971), .B2(n387), .ZN(n2408)
         );
  OAI22_X2 U2056 ( .A1(n3416), .A2(n2973), .B1(n2972), .B2(n387), .ZN(n2409)
         );
  OAI22_X2 U2057 ( .A1(n3416), .A2(n2974), .B1(n2973), .B2(n387), .ZN(n2410)
         );
  OAI22_X2 U2058 ( .A1(n3416), .A2(n2975), .B1(n2974), .B2(n387), .ZN(n2411)
         );
  OAI22_X2 U2060 ( .A1(n3416), .A2(n2977), .B1(n2976), .B2(n387), .ZN(n2413)
         );
  OAI22_X2 U2062 ( .A1(n3416), .A2(n2979), .B1(n2978), .B2(n387), .ZN(n2415)
         );
  OAI22_X2 U2063 ( .A1(n3416), .A2(n2980), .B1(n2979), .B2(n387), .ZN(n2416)
         );
  OAI22_X2 U2064 ( .A1(n3416), .A2(n2981), .B1(n2980), .B2(n387), .ZN(n2417)
         );
  OAI22_X2 U2066 ( .A1(n3416), .A2(n2983), .B1(n2982), .B2(n387), .ZN(n2419)
         );
  OAI22_X2 U2067 ( .A1(n3416), .A2(n2984), .B1(n2983), .B2(n387), .ZN(n2420)
         );
  OAI22_X2 U2068 ( .A1(n3416), .A2(n2985), .B1(n2984), .B2(n387), .ZN(n2421)
         );
  OAI22_X2 U2069 ( .A1(n3416), .A2(n2986), .B1(n2985), .B2(n387), .ZN(n2422)
         );
  OAI22_X2 U2070 ( .A1(n3416), .A2(n2987), .B1(n2986), .B2(n387), .ZN(n2423)
         );
  OAI22_X2 U2071 ( .A1(n3416), .A2(n2988), .B1(n2987), .B2(n387), .ZN(n2424)
         );
  OAI22_X2 U2072 ( .A1(n3416), .A2(n2989), .B1(n2988), .B2(n387), .ZN(n2425)
         );
  OAI22_X2 U2073 ( .A1(n3416), .A2(n2990), .B1(n2989), .B2(n387), .ZN(n2426)
         );
  OAI22_X2 U2074 ( .A1(n3416), .A2(n2991), .B1(n2990), .B2(n387), .ZN(n2427)
         );
  OAI22_X2 U2075 ( .A1(n3416), .A2(n2992), .B1(n2991), .B2(n387), .ZN(n2428)
         );
  OAI22_X2 U2076 ( .A1(n3416), .A2(n2993), .B1(n2992), .B2(n387), .ZN(n2429)
         );
  OAI22_X2 U2077 ( .A1(n3416), .A2(n2994), .B1(n2993), .B2(n387), .ZN(n2430)
         );
  OAI22_X2 U2078 ( .A1(n3416), .A2(n2995), .B1(n2994), .B2(n387), .ZN(n2431)
         );
  OAI22_X2 U2079 ( .A1(n3416), .A2(n2996), .B1(n2995), .B2(n387), .ZN(n2432)
         );
  OAI22_X2 U2112 ( .A1(n434), .A2(n3287), .B1(n3030), .B2(n3641), .ZN(n2071)
         );
  OAI22_X2 U2113 ( .A1(n434), .A2(n2998), .B1(n3641), .B2(n3287), .ZN(n2435)
         );
  OAI22_X2 U2116 ( .A1(n434), .A2(n3001), .B1(n3000), .B2(n3641), .ZN(n2438)
         );
  OAI22_X2 U2119 ( .A1(n434), .A2(n3004), .B1(n3003), .B2(n3641), .ZN(n2441)
         );
  OAI22_X2 U2123 ( .A1(n434), .A2(n3008), .B1(n3007), .B2(n3641), .ZN(n2445)
         );
  OAI22_X2 U2124 ( .A1(n434), .A2(n3009), .B1(n3008), .B2(n3641), .ZN(n2446)
         );
  OAI22_X2 U2125 ( .A1(n434), .A2(n3010), .B1(n3009), .B2(n3641), .ZN(n2447)
         );
  OAI22_X2 U2126 ( .A1(n434), .A2(n3011), .B1(n3010), .B2(n3641), .ZN(n2448)
         );
  OAI22_X2 U2132 ( .A1(n434), .A2(n3017), .B1(n3016), .B2(n3641), .ZN(n2454)
         );
  OAI22_X2 U2133 ( .A1(n434), .A2(n3018), .B1(n3017), .B2(n3641), .ZN(n2455)
         );
  OAI22_X2 U2135 ( .A1(n434), .A2(n3020), .B1(n3019), .B2(n3641), .ZN(n2457)
         );
  OAI22_X2 U2136 ( .A1(n434), .A2(n3021), .B1(n3020), .B2(n3641), .ZN(n2458)
         );
  OAI22_X2 U2140 ( .A1(n434), .A2(n3025), .B1(n3024), .B2(n3641), .ZN(n2462)
         );
  OAI22_X2 U2143 ( .A1(n434), .A2(n3028), .B1(n3027), .B2(n3641), .ZN(n2465)
         );
  OAI22_X2 U2144 ( .A1(n434), .A2(n3029), .B1(n3028), .B2(n3641), .ZN(n2466)
         );
  OAI22_X2 U2181 ( .A1(n3560), .A2(n3034), .B1(n3033), .B2(n381), .ZN(n2472)
         );
  OAI22_X2 U2183 ( .A1(n3560), .A2(n3036), .B1(n3035), .B2(n381), .ZN(n2474)
         );
  OAI22_X2 U2185 ( .A1(n3560), .A2(n3038), .B1(n3037), .B2(n381), .ZN(n2476)
         );
  OAI22_X2 U2202 ( .A1(n3560), .A2(n3055), .B1(n3054), .B2(n381), .ZN(n2493)
         );
  OAI22_X2 U2204 ( .A1(n3560), .A2(n3057), .B1(n3056), .B2(n381), .ZN(n2495)
         );
  OAI22_X2 U2372 ( .A1(n3555), .A2(n3291), .B1(n3162), .B2(n372), .ZN(n2075)
         );
  OAI22_X2 U2373 ( .A1(n422), .A2(n3130), .B1(n372), .B2(n3291), .ZN(n2571) );
  OAI22_X2 U2376 ( .A1(n422), .A2(n3133), .B1(n3132), .B2(n372), .ZN(n2574) );
  OAI22_X2 U2377 ( .A1(n422), .A2(n3134), .B1(n3133), .B2(n372), .ZN(n2575) );
  OAI22_X2 U2378 ( .A1(n422), .A2(n3135), .B1(n3134), .B2(n372), .ZN(n2576) );
  OAI22_X2 U2379 ( .A1(n422), .A2(n3136), .B1(n3135), .B2(n372), .ZN(n2577) );
  OAI22_X2 U2380 ( .A1(n422), .A2(n3137), .B1(n3136), .B2(n372), .ZN(n2578) );
  OAI22_X2 U2381 ( .A1(n422), .A2(n3138), .B1(n3137), .B2(n372), .ZN(n2579) );
  OAI22_X2 U2382 ( .A1(n422), .A2(n3139), .B1(n3138), .B2(n372), .ZN(n2580) );
  OAI22_X2 U2383 ( .A1(n422), .A2(n3140), .B1(n3139), .B2(n372), .ZN(n2581) );
  OAI22_X2 U2384 ( .A1(n422), .A2(n3141), .B1(n3140), .B2(n372), .ZN(n2582) );
  OAI22_X2 U2385 ( .A1(n422), .A2(n3142), .B1(n3141), .B2(n372), .ZN(n2583) );
  OAI22_X2 U2387 ( .A1(n422), .A2(n3144), .B1(n3143), .B2(n372), .ZN(n2585) );
  OAI22_X2 U2388 ( .A1(n422), .A2(n3145), .B1(n3144), .B2(n372), .ZN(n2586) );
  OAI22_X2 U2389 ( .A1(n422), .A2(n3146), .B1(n3145), .B2(n372), .ZN(n2587) );
  OAI22_X2 U2390 ( .A1(n3555), .A2(n3147), .B1(n3146), .B2(n372), .ZN(n2588)
         );
  OAI22_X2 U2391 ( .A1(n422), .A2(n3148), .B1(n3147), .B2(n372), .ZN(n2589) );
  OAI22_X2 U2392 ( .A1(n422), .A2(n3149), .B1(n3148), .B2(n372), .ZN(n2590) );
  OAI22_X2 U2393 ( .A1(n422), .A2(n3150), .B1(n3149), .B2(n372), .ZN(n2591) );
  OAI22_X2 U2394 ( .A1(n422), .A2(n3151), .B1(n3150), .B2(n372), .ZN(n2592) );
  OAI22_X2 U2395 ( .A1(n422), .A2(n3152), .B1(n3151), .B2(n372), .ZN(n2593) );
  OAI22_X2 U2396 ( .A1(n422), .A2(n3153), .B1(n3152), .B2(n372), .ZN(n2594) );
  OAI22_X2 U2397 ( .A1(n422), .A2(n3154), .B1(n3153), .B2(n372), .ZN(n2595) );
  OAI22_X2 U2398 ( .A1(n422), .A2(n3155), .B1(n3154), .B2(n372), .ZN(n2596) );
  OAI22_X2 U2399 ( .A1(n422), .A2(n3156), .B1(n3155), .B2(n372), .ZN(n2597) );
  OAI22_X2 U2400 ( .A1(n422), .A2(n3157), .B1(n3156), .B2(n372), .ZN(n2598) );
  OAI22_X2 U2401 ( .A1(n3555), .A2(n3158), .B1(n3157), .B2(n372), .ZN(n2599)
         );
  OAI22_X2 U2402 ( .A1(n3555), .A2(n3159), .B1(n3158), .B2(n372), .ZN(n2600)
         );
  OAI22_X2 U2403 ( .A1(n3555), .A2(n3160), .B1(n3159), .B2(n372), .ZN(n2601)
         );
  OAI22_X2 U2404 ( .A1(n422), .A2(n3161), .B1(n3160), .B2(n372), .ZN(n2602) );
  OAI22_X2 U2439 ( .A1(n419), .A2(n3164), .B1(n3163), .B2(n369), .ZN(n2606) );
  OAI22_X2 U2440 ( .A1(n419), .A2(n3165), .B1(n3164), .B2(n369), .ZN(n2607) );
  OAI22_X2 U2441 ( .A1(n419), .A2(n3166), .B1(n3165), .B2(n369), .ZN(n2608) );
  OAI22_X2 U2442 ( .A1(n419), .A2(n3167), .B1(n3166), .B2(n369), .ZN(n2609) );
  OAI22_X2 U2443 ( .A1(n419), .A2(n3168), .B1(n3167), .B2(n369), .ZN(n2610) );
  OAI22_X2 U2444 ( .A1(n419), .A2(n3169), .B1(n3168), .B2(n369), .ZN(n2611) );
  OAI22_X2 U2445 ( .A1(n419), .A2(n3170), .B1(n3169), .B2(n369), .ZN(n2612) );
  OAI22_X2 U2446 ( .A1(n419), .A2(n3171), .B1(n3170), .B2(n369), .ZN(n2613) );
  OAI22_X2 U2447 ( .A1(n419), .A2(n3172), .B1(n3171), .B2(n369), .ZN(n2614) );
  OAI22_X2 U2448 ( .A1(n419), .A2(n3173), .B1(n3172), .B2(n369), .ZN(n2615) );
  OAI22_X2 U2449 ( .A1(n419), .A2(n3174), .B1(n3173), .B2(n369), .ZN(n2616) );
  OAI22_X2 U2450 ( .A1(n419), .A2(n3175), .B1(n3174), .B2(n369), .ZN(n2617) );
  OAI22_X2 U2451 ( .A1(n419), .A2(n3176), .B1(n3175), .B2(n369), .ZN(n2618) );
  OAI22_X2 U2452 ( .A1(n419), .A2(n3177), .B1(n3176), .B2(n369), .ZN(n2619) );
  OAI22_X2 U2453 ( .A1(n419), .A2(n3178), .B1(n3177), .B2(n369), .ZN(n2620) );
  OAI22_X2 U2454 ( .A1(n419), .A2(n3179), .B1(n3178), .B2(n369), .ZN(n2621) );
  OAI22_X2 U2455 ( .A1(n419), .A2(n3180), .B1(n3179), .B2(n369), .ZN(n2622) );
  OAI22_X2 U2456 ( .A1(n419), .A2(n3181), .B1(n3180), .B2(n369), .ZN(n2623) );
  OAI22_X2 U2457 ( .A1(n419), .A2(n3182), .B1(n3181), .B2(n369), .ZN(n2624) );
  OAI22_X2 U2458 ( .A1(n419), .A2(n3183), .B1(n3182), .B2(n369), .ZN(n2625) );
  OAI22_X2 U2459 ( .A1(n419), .A2(n3184), .B1(n3183), .B2(n369), .ZN(n2626) );
  OAI22_X2 U2460 ( .A1(n419), .A2(n3185), .B1(n3184), .B2(n369), .ZN(n2627) );
  OAI22_X2 U2461 ( .A1(n419), .A2(n3186), .B1(n3185), .B2(n369), .ZN(n2628) );
  OAI22_X2 U2462 ( .A1(n419), .A2(n3187), .B1(n3186), .B2(n369), .ZN(n2629) );
  OAI22_X2 U2463 ( .A1(n419), .A2(n3188), .B1(n3187), .B2(n369), .ZN(n2630) );
  OAI22_X2 U2464 ( .A1(n419), .A2(n3189), .B1(n3188), .B2(n369), .ZN(n2631) );
  OAI22_X2 U2465 ( .A1(n419), .A2(n3190), .B1(n3189), .B2(n369), .ZN(n2632) );
  OAI22_X2 U2466 ( .A1(n419), .A2(n3191), .B1(n3190), .B2(n369), .ZN(n2633) );
  OAI22_X2 U2467 ( .A1(n419), .A2(n3192), .B1(n3191), .B2(n369), .ZN(n2634) );
  OAI22_X2 U2468 ( .A1(n419), .A2(n3193), .B1(n3192), .B2(n369), .ZN(n2635) );
  OAI22_X2 U2469 ( .A1(n419), .A2(n3194), .B1(n3193), .B2(n369), .ZN(n2636) );
  XOR2_X2 U2548 ( .A(n354), .B(a[22]), .Z(n3232) );
  XOR2_X2 U2554 ( .A(n3425), .B(n348), .Z(n3234) );
  XOR2_X2 U2572 ( .A(a[6]), .B(n330), .Z(n3240) );
  INV_X4 U2585 ( .A(a[16]), .ZN(n3781) );
  INV_X2 U2586 ( .A(a[26]), .ZN(n3755) );
  INV_X2 U2587 ( .A(n3501), .ZN(n3502) );
  INV_X2 U2588 ( .A(n3563), .ZN(n3556) );
  INV_X1 U2589 ( .A(n351), .ZN(n3585) );
  INV_X1 U2590 ( .A(n342), .ZN(n3633) );
  INV_X1 U2591 ( .A(n342), .ZN(n3608) );
  INV_X2 U2592 ( .A(n348), .ZN(n3644) );
  INV_X1 U2593 ( .A(n366), .ZN(n416) );
  INV_X2 U2594 ( .A(n330), .ZN(n3667) );
  INV_X1 U2595 ( .A(n363), .ZN(n3278) );
  INV_X1 U2596 ( .A(n363), .ZN(n3482) );
  BUF_X1 U2597 ( .A(n357), .Z(n3467) );
  XNOR2_X1 U2598 ( .A(n3781), .B(n345), .ZN(n3235) );
  INV_X2 U2599 ( .A(n345), .ZN(n3563) );
  XNOR2_X1 U2600 ( .A(n465), .B(n321), .ZN(n3194) );
  XNOR2_X1 U2601 ( .A(n465), .B(n327), .ZN(n3128) );
  XNOR2_X1 U2602 ( .A(n465), .B(n333), .ZN(n3062) );
  XNOR2_X1 U2603 ( .A(n465), .B(n3778), .ZN(n3161) );
  XNOR2_X1 U2604 ( .A(n465), .B(n336), .ZN(n3029) );
  XNOR2_X1 U2605 ( .A(n465), .B(n3564), .ZN(n2930) );
  AND2_X1 U2606 ( .A1(n465), .A2(n366), .ZN(n2093) );
  XNOR2_X1 U2607 ( .A(n465), .B(n351), .ZN(n2864) );
  XNOR2_X1 U2608 ( .A(n465), .B(n360), .ZN(n2765) );
  XNOR2_X1 U2609 ( .A(n465), .B(n354), .ZN(n2831) );
  XNOR2_X1 U2610 ( .A(n465), .B(n339), .ZN(n2996) );
  XNOR2_X1 U2611 ( .A(n465), .B(n3634), .ZN(n2963) );
  XNOR2_X1 U2612 ( .A(n465), .B(n3645), .ZN(n2897) );
  XNOR2_X1 U2613 ( .A(n465), .B(n330), .ZN(n3095) );
  XNOR2_X1 U2614 ( .A(n465), .B(n366), .ZN(n2699) );
  XNOR2_X1 U2615 ( .A(n465), .B(n363), .ZN(n2732) );
  XNOR2_X1 U2616 ( .A(n465), .B(n357), .ZN(n2798) );
  INV_X2 U2617 ( .A(a[10]), .ZN(n3752) );
  INV_X2 U2618 ( .A(a[2]), .ZN(n3737) );
  INV_X2 U2619 ( .A(a[12]), .ZN(n3758) );
  INV_X2 U2620 ( .A(a[20]), .ZN(n3760) );
  INV_X2 U2621 ( .A(a[8]), .ZN(n3767) );
  XOR2_X1 U2622 ( .A(a[14]), .B(n342), .Z(n3236) );
  INV_X2 U2623 ( .A(a[14]), .ZN(n3762) );
  INV_X2 U2624 ( .A(a[22]), .ZN(n3629) );
  AND2_X1 U2625 ( .A1(n465), .A2(a[0]), .ZN(product[0]) );
  OAI21_X1 U2626 ( .B1(a[0]), .B2(n3785), .A(n321), .ZN(n2604) );
  XNOR2_X1 U2627 ( .A(a[0]), .B(n321), .ZN(n3529) );
  XNOR2_X1 U2628 ( .A(n3737), .B(n324), .ZN(n3242) );
  INV_X2 U2629 ( .A(n324), .ZN(n3777) );
  INV_X1 U2630 ( .A(n324), .ZN(n3501) );
  INV_X1 U2631 ( .A(n511), .ZN(n2646) );
  XNOR2_X1 U2632 ( .A(n511), .B(n360), .ZN(n2743) );
  XNOR2_X1 U2633 ( .A(n511), .B(n363), .ZN(n2710) );
  XNOR2_X1 U2634 ( .A(n511), .B(n3645), .ZN(n2875) );
  XNOR2_X1 U2635 ( .A(n511), .B(n366), .ZN(n2677) );
  XNOR2_X1 U2636 ( .A(n511), .B(n321), .ZN(n3172) );
  XNOR2_X1 U2637 ( .A(n511), .B(n339), .ZN(n2974) );
  XNOR2_X1 U2638 ( .A(n511), .B(n351), .ZN(n2842) );
  XNOR2_X1 U2639 ( .A(n511), .B(n330), .ZN(n3073) );
  XNOR2_X1 U2640 ( .A(n511), .B(n336), .ZN(n3007) );
  XNOR2_X1 U2641 ( .A(n511), .B(n357), .ZN(n2776) );
  XNOR2_X1 U2642 ( .A(n511), .B(n3502), .ZN(n3139) );
  XNOR2_X1 U2643 ( .A(n511), .B(n342), .ZN(n2941) );
  XNOR2_X1 U2644 ( .A(n511), .B(n354), .ZN(n2809) );
  XNOR2_X1 U2645 ( .A(n511), .B(n333), .ZN(n3040) );
  XNOR2_X1 U2646 ( .A(n511), .B(n345), .ZN(n2908) );
  INV_X1 U2647 ( .A(n505), .ZN(n2649) );
  XNOR2_X1 U2648 ( .A(n505), .B(n366), .ZN(n2680) );
  XNOR2_X1 U2649 ( .A(n505), .B(n336), .ZN(n3010) );
  XNOR2_X1 U2650 ( .A(n505), .B(n342), .ZN(n2944) );
  XNOR2_X1 U2651 ( .A(n505), .B(n363), .ZN(n2713) );
  XNOR2_X1 U2652 ( .A(n505), .B(n348), .ZN(n2878) );
  XNOR2_X1 U2653 ( .A(n505), .B(n351), .ZN(n2845) );
  XNOR2_X1 U2654 ( .A(n505), .B(n354), .ZN(n2812) );
  XNOR2_X1 U2655 ( .A(n505), .B(n360), .ZN(n2746) );
  XNOR2_X1 U2656 ( .A(n505), .B(n357), .ZN(n2779) );
  XNOR2_X1 U2657 ( .A(n505), .B(n327), .ZN(n3109) );
  XNOR2_X1 U2658 ( .A(n505), .B(n339), .ZN(n2977) );
  XNOR2_X1 U2659 ( .A(n505), .B(n321), .ZN(n3175) );
  XNOR2_X1 U2660 ( .A(n505), .B(n345), .ZN(n2911) );
  XNOR2_X1 U2661 ( .A(n505), .B(n324), .ZN(n3142) );
  XNOR2_X1 U2662 ( .A(n505), .B(n333), .ZN(n3043) );
  XNOR2_X1 U2663 ( .A(n505), .B(n330), .ZN(n3076) );
  INV_X1 U2664 ( .A(n513), .ZN(n2645) );
  XNOR2_X1 U2665 ( .A(n513), .B(n360), .ZN(n2742) );
  XNOR2_X1 U2666 ( .A(n513), .B(n363), .ZN(n2709) );
  XNOR2_X1 U2667 ( .A(n513), .B(n354), .ZN(n2808) );
  XNOR2_X1 U2668 ( .A(n513), .B(n342), .ZN(n2940) );
  XNOR2_X1 U2669 ( .A(n513), .B(n366), .ZN(n2676) );
  XNOR2_X1 U2670 ( .A(n513), .B(n351), .ZN(n2841) );
  XNOR2_X1 U2671 ( .A(n513), .B(n348), .ZN(n2874) );
  XNOR2_X1 U2672 ( .A(n513), .B(n336), .ZN(n3006) );
  XNOR2_X1 U2673 ( .A(n513), .B(n339), .ZN(n2973) );
  XNOR2_X1 U2674 ( .A(n513), .B(n333), .ZN(n3039) );
  XNOR2_X1 U2675 ( .A(n513), .B(n321), .ZN(n3171) );
  XNOR2_X1 U2676 ( .A(n513), .B(n357), .ZN(n2775) );
  XNOR2_X1 U2677 ( .A(n513), .B(n324), .ZN(n3138) );
  XNOR2_X1 U2678 ( .A(n513), .B(n330), .ZN(n3072) );
  XNOR2_X1 U2679 ( .A(n513), .B(n327), .ZN(n3105) );
  XNOR2_X1 U2680 ( .A(n513), .B(n345), .ZN(n2907) );
  INV_X1 U2681 ( .A(n499), .ZN(n2652) );
  XNOR2_X1 U2682 ( .A(n499), .B(n366), .ZN(n2683) );
  XNOR2_X1 U2683 ( .A(n499), .B(n3467), .ZN(n2782) );
  XNOR2_X1 U2684 ( .A(n499), .B(n360), .ZN(n2749) );
  XNOR2_X1 U2685 ( .A(n499), .B(n330), .ZN(n3079) );
  XNOR2_X1 U2686 ( .A(n499), .B(n363), .ZN(n2716) );
  XNOR2_X1 U2687 ( .A(n499), .B(n339), .ZN(n2980) );
  XNOR2_X1 U2688 ( .A(n499), .B(n327), .ZN(n3112) );
  XNOR2_X1 U2689 ( .A(n499), .B(n348), .ZN(n2881) );
  XNOR2_X1 U2690 ( .A(n499), .B(n3556), .ZN(n2914) );
  XNOR2_X1 U2691 ( .A(n499), .B(n324), .ZN(n3145) );
  XNOR2_X1 U2692 ( .A(n499), .B(n321), .ZN(n3178) );
  XNOR2_X1 U2693 ( .A(n499), .B(n342), .ZN(n2947) );
  XNOR2_X1 U2694 ( .A(n499), .B(n336), .ZN(n3013) );
  XNOR2_X1 U2695 ( .A(n499), .B(n333), .ZN(n3046) );
  XNOR2_X1 U2696 ( .A(n499), .B(n354), .ZN(n2815) );
  XNOR2_X1 U2697 ( .A(n499), .B(n351), .ZN(n2848) );
  INV_X1 U2698 ( .A(n507), .ZN(n2648) );
  XNOR2_X1 U2699 ( .A(n507), .B(n363), .ZN(n2712) );
  XNOR2_X1 U2700 ( .A(n507), .B(n366), .ZN(n2679) );
  XNOR2_X1 U2701 ( .A(n507), .B(n342), .ZN(n2943) );
  XNOR2_X1 U2702 ( .A(n507), .B(n333), .ZN(n3042) );
  XNOR2_X1 U2703 ( .A(n507), .B(n351), .ZN(n2844) );
  XNOR2_X1 U2704 ( .A(n507), .B(n3502), .ZN(n3141) );
  XNOR2_X1 U2705 ( .A(n507), .B(n360), .ZN(n2745) );
  XNOR2_X1 U2706 ( .A(n507), .B(n354), .ZN(n2811) );
  XNOR2_X1 U2707 ( .A(n507), .B(n357), .ZN(n2778) );
  XNOR2_X1 U2708 ( .A(n507), .B(n336), .ZN(n3009) );
  XNOR2_X1 U2709 ( .A(n507), .B(n330), .ZN(n3075) );
  XNOR2_X1 U2710 ( .A(n507), .B(n327), .ZN(n3108) );
  XNOR2_X1 U2711 ( .A(n507), .B(n339), .ZN(n2976) );
  XNOR2_X1 U2712 ( .A(n507), .B(n345), .ZN(n2910) );
  XNOR2_X1 U2713 ( .A(n507), .B(n321), .ZN(n3174) );
  INV_X1 U2714 ( .A(n501), .ZN(n2651) );
  XNOR2_X1 U2715 ( .A(n501), .B(n366), .ZN(n2682) );
  XNOR2_X1 U2716 ( .A(n501), .B(n3467), .ZN(n2781) );
  XNOR2_X1 U2717 ( .A(n501), .B(n327), .ZN(n3111) );
  XNOR2_X1 U2718 ( .A(n501), .B(n363), .ZN(n2715) );
  XNOR2_X1 U2719 ( .A(n501), .B(n330), .ZN(n3078) );
  XNOR2_X1 U2720 ( .A(n501), .B(n3564), .ZN(n2913) );
  XNOR2_X1 U2721 ( .A(n501), .B(n360), .ZN(n2748) );
  XNOR2_X1 U2722 ( .A(n501), .B(n324), .ZN(n3144) );
  XNOR2_X1 U2723 ( .A(n501), .B(n348), .ZN(n2880) );
  XNOR2_X1 U2724 ( .A(n501), .B(n339), .ZN(n2979) );
  XNOR2_X1 U2725 ( .A(n501), .B(n342), .ZN(n2946) );
  XNOR2_X1 U2726 ( .A(n501), .B(n336), .ZN(n3012) );
  XNOR2_X1 U2727 ( .A(n501), .B(n333), .ZN(n3045) );
  XNOR2_X1 U2728 ( .A(n501), .B(n321), .ZN(n3177) );
  XNOR2_X1 U2729 ( .A(n501), .B(n354), .ZN(n2814) );
  XNOR2_X1 U2730 ( .A(n501), .B(n351), .ZN(n2847) );
  INV_X1 U2731 ( .A(n493), .ZN(n2655) );
  XNOR2_X1 U2732 ( .A(n493), .B(n351), .ZN(n2851) );
  XNOR2_X1 U2733 ( .A(n493), .B(n333), .ZN(n3049) );
  XNOR2_X1 U2734 ( .A(n493), .B(n363), .ZN(n2719) );
  XNOR2_X1 U2735 ( .A(n493), .B(n336), .ZN(n3016) );
  XNOR2_X1 U2736 ( .A(n493), .B(n342), .ZN(n2950) );
  XNOR2_X1 U2737 ( .A(n493), .B(n360), .ZN(n2752) );
  XNOR2_X1 U2738 ( .A(n493), .B(n348), .ZN(n2884) );
  XNOR2_X1 U2739 ( .A(n493), .B(n345), .ZN(n2917) );
  XNOR2_X1 U2740 ( .A(n493), .B(n330), .ZN(n3082) );
  XNOR2_X1 U2741 ( .A(n493), .B(n366), .ZN(n2686) );
  XNOR2_X1 U2742 ( .A(n493), .B(n321), .ZN(n3181) );
  XNOR2_X1 U2743 ( .A(n493), .B(n354), .ZN(n2818) );
  XNOR2_X1 U2744 ( .A(n493), .B(n327), .ZN(n3115) );
  XNOR2_X1 U2745 ( .A(n493), .B(n357), .ZN(n2785) );
  XNOR2_X1 U2746 ( .A(n493), .B(n3502), .ZN(n3148) );
  XNOR2_X1 U2747 ( .A(n493), .B(n339), .ZN(n2983) );
  INV_X1 U2748 ( .A(n495), .ZN(n2654) );
  XNOR2_X1 U2749 ( .A(n495), .B(n351), .ZN(n2850) );
  XNOR2_X1 U2750 ( .A(n495), .B(n333), .ZN(n3048) );
  XNOR2_X1 U2751 ( .A(n495), .B(n360), .ZN(n2751) );
  XNOR2_X1 U2752 ( .A(n495), .B(n366), .ZN(n2685) );
  XNOR2_X1 U2753 ( .A(n495), .B(n363), .ZN(n2718) );
  XNOR2_X1 U2754 ( .A(n495), .B(n3556), .ZN(n2916) );
  XNOR2_X1 U2755 ( .A(n495), .B(n3502), .ZN(n3147) );
  XNOR2_X1 U2756 ( .A(n495), .B(n348), .ZN(n2883) );
  XNOR2_X1 U2757 ( .A(n495), .B(n336), .ZN(n3015) );
  XNOR2_X1 U2758 ( .A(n495), .B(n330), .ZN(n3081) );
  XNOR2_X1 U2759 ( .A(n495), .B(n342), .ZN(n2949) );
  XNOR2_X1 U2760 ( .A(n495), .B(n357), .ZN(n2784) );
  XNOR2_X1 U2761 ( .A(n495), .B(n354), .ZN(n2817) );
  XNOR2_X1 U2762 ( .A(n495), .B(n339), .ZN(n2982) );
  XNOR2_X1 U2763 ( .A(n495), .B(n327), .ZN(n3114) );
  XNOR2_X1 U2764 ( .A(n495), .B(n321), .ZN(n3180) );
  INV_X1 U2765 ( .A(n489), .ZN(n2657) );
  XNOR2_X1 U2766 ( .A(n489), .B(n333), .ZN(n3051) );
  XNOR2_X1 U2767 ( .A(n489), .B(n330), .ZN(n3084) );
  XNOR2_X1 U2768 ( .A(n489), .B(n366), .ZN(n2688) );
  XNOR2_X1 U2769 ( .A(n489), .B(n363), .ZN(n2721) );
  XNOR2_X1 U2770 ( .A(n489), .B(n354), .ZN(n2820) );
  XNOR2_X1 U2771 ( .A(n489), .B(n321), .ZN(n3183) );
  XNOR2_X1 U2772 ( .A(n489), .B(n327), .ZN(n3117) );
  XNOR2_X1 U2773 ( .A(n489), .B(n348), .ZN(n2886) );
  XNOR2_X1 U2774 ( .A(n489), .B(n339), .ZN(n2985) );
  XNOR2_X1 U2775 ( .A(n489), .B(n336), .ZN(n3018) );
  XNOR2_X1 U2776 ( .A(n489), .B(n342), .ZN(n2952) );
  XNOR2_X1 U2777 ( .A(n489), .B(n351), .ZN(n2853) );
  XNOR2_X1 U2778 ( .A(n489), .B(n3556), .ZN(n2919) );
  XNOR2_X1 U2779 ( .A(n489), .B(n360), .ZN(n2754) );
  XNOR2_X1 U2780 ( .A(n489), .B(n3502), .ZN(n3150) );
  INV_X1 U2781 ( .A(n483), .ZN(n2660) );
  XNOR2_X1 U2782 ( .A(n483), .B(n342), .ZN(n2955) );
  XNOR2_X1 U2783 ( .A(n483), .B(n321), .ZN(n3186) );
  XNOR2_X1 U2784 ( .A(n483), .B(n366), .ZN(n2691) );
  XNOR2_X1 U2785 ( .A(n483), .B(n363), .ZN(n2724) );
  XNOR2_X1 U2786 ( .A(n483), .B(n327), .ZN(n3120) );
  XNOR2_X1 U2787 ( .A(n483), .B(n354), .ZN(n2823) );
  XNOR2_X1 U2788 ( .A(n483), .B(n333), .ZN(n3054) );
  XNOR2_X1 U2789 ( .A(n483), .B(n3513), .ZN(n3153) );
  XNOR2_X1 U2790 ( .A(n483), .B(n348), .ZN(n2889) );
  XNOR2_X1 U2791 ( .A(n483), .B(n351), .ZN(n2856) );
  XNOR2_X1 U2792 ( .A(n483), .B(n330), .ZN(n3087) );
  XNOR2_X1 U2793 ( .A(n483), .B(n339), .ZN(n2988) );
  XNOR2_X1 U2794 ( .A(n483), .B(n360), .ZN(n2757) );
  XNOR2_X1 U2795 ( .A(n483), .B(n357), .ZN(n2790) );
  XNOR2_X1 U2796 ( .A(n483), .B(n3556), .ZN(n2922) );
  XNOR2_X1 U2797 ( .A(n483), .B(n336), .ZN(n3021) );
  XNOR2_X1 U2798 ( .A(n477), .B(n330), .ZN(n3090) );
  INV_X1 U2799 ( .A(n477), .ZN(n2663) );
  XNOR2_X1 U2800 ( .A(n477), .B(n321), .ZN(n3189) );
  XNOR2_X1 U2801 ( .A(n477), .B(n3513), .ZN(n3156) );
  XNOR2_X1 U2802 ( .A(n477), .B(n3634), .ZN(n2958) );
  XNOR2_X1 U2803 ( .A(n477), .B(n327), .ZN(n3123) );
  XNOR2_X1 U2804 ( .A(n477), .B(n354), .ZN(n2826) );
  XNOR2_X1 U2805 ( .A(n477), .B(n348), .ZN(n2892) );
  XNOR2_X1 U2806 ( .A(n477), .B(n336), .ZN(n3024) );
  XNOR2_X1 U2807 ( .A(n477), .B(n357), .ZN(n2793) );
  XNOR2_X1 U2808 ( .A(n477), .B(n339), .ZN(n2991) );
  XNOR2_X1 U2809 ( .A(n477), .B(n366), .ZN(n2694) );
  XNOR2_X1 U2810 ( .A(n477), .B(n333), .ZN(n3057) );
  XNOR2_X1 U2811 ( .A(n477), .B(n360), .ZN(n2760) );
  XNOR2_X1 U2812 ( .A(n477), .B(n3556), .ZN(n2925) );
  XNOR2_X1 U2813 ( .A(n477), .B(n363), .ZN(n2727) );
  XNOR2_X1 U2814 ( .A(n477), .B(n351), .ZN(n2859) );
  INV_X1 U2815 ( .A(n487), .ZN(n2658) );
  XNOR2_X1 U2816 ( .A(n487), .B(n363), .ZN(n2722) );
  XNOR2_X1 U2817 ( .A(n487), .B(n366), .ZN(n2689) );
  XNOR2_X1 U2818 ( .A(n487), .B(n330), .ZN(n3085) );
  XNOR2_X1 U2819 ( .A(n487), .B(n327), .ZN(n3118) );
  XNOR2_X1 U2820 ( .A(n487), .B(n321), .ZN(n3184) );
  XNOR2_X1 U2821 ( .A(n487), .B(n339), .ZN(n2986) );
  XNOR2_X1 U2822 ( .A(n487), .B(n3513), .ZN(n3151) );
  XNOR2_X1 U2823 ( .A(n487), .B(n336), .ZN(n3019) );
  XNOR2_X1 U2824 ( .A(n487), .B(n351), .ZN(n2854) );
  XNOR2_X1 U2825 ( .A(n487), .B(n354), .ZN(n2821) );
  XNOR2_X1 U2826 ( .A(n487), .B(n342), .ZN(n2953) );
  XNOR2_X1 U2827 ( .A(n487), .B(n360), .ZN(n2755) );
  XNOR2_X1 U2828 ( .A(n487), .B(n333), .ZN(n3052) );
  INV_X1 U2829 ( .A(n481), .ZN(n2661) );
  XNOR2_X1 U2830 ( .A(n481), .B(n321), .ZN(n3187) );
  XNOR2_X1 U2831 ( .A(n481), .B(n351), .ZN(n2857) );
  XNOR2_X1 U2832 ( .A(n481), .B(n3513), .ZN(n3154) );
  XNOR2_X1 U2833 ( .A(n481), .B(n330), .ZN(n3088) );
  XNOR2_X1 U2834 ( .A(n481), .B(n333), .ZN(n3055) );
  XNOR2_X1 U2835 ( .A(n481), .B(n354), .ZN(n2824) );
  XNOR2_X1 U2836 ( .A(n481), .B(n339), .ZN(n2989) );
  XNOR2_X1 U2837 ( .A(n481), .B(n327), .ZN(n3121) );
  XNOR2_X1 U2838 ( .A(n481), .B(n366), .ZN(n2692) );
  XNOR2_X1 U2839 ( .A(n481), .B(n363), .ZN(n2725) );
  XNOR2_X1 U2840 ( .A(n481), .B(n360), .ZN(n2758) );
  XNOR2_X1 U2841 ( .A(n481), .B(n342), .ZN(n2956) );
  XNOR2_X1 U2842 ( .A(n481), .B(n3564), .ZN(n2923) );
  XNOR2_X1 U2843 ( .A(n481), .B(n336), .ZN(n3022) );
  XNOR2_X1 U2844 ( .A(n481), .B(n348), .ZN(n2890) );
  XNOR2_X1 U2845 ( .A(n481), .B(n357), .ZN(n2791) );
  XNOR2_X1 U2846 ( .A(n475), .B(n321), .ZN(n3190) );
  XNOR2_X1 U2847 ( .A(n475), .B(n3513), .ZN(n3157) );
  XNOR2_X1 U2848 ( .A(n475), .B(n327), .ZN(n3124) );
  INV_X1 U2849 ( .A(n475), .ZN(n2664) );
  XNOR2_X1 U2850 ( .A(n475), .B(n333), .ZN(n3058) );
  XNOR2_X1 U2851 ( .A(n475), .B(n348), .ZN(n2893) );
  XNOR2_X1 U2852 ( .A(n475), .B(n330), .ZN(n3091) );
  XNOR2_X1 U2853 ( .A(n475), .B(n354), .ZN(n2827) );
  XNOR2_X1 U2854 ( .A(n475), .B(n366), .ZN(n2695) );
  XNOR2_X1 U2855 ( .A(n475), .B(n339), .ZN(n2992) );
  XNOR2_X1 U2856 ( .A(n475), .B(n342), .ZN(n2959) );
  XNOR2_X1 U2857 ( .A(n475), .B(n360), .ZN(n2761) );
  XNOR2_X1 U2858 ( .A(n475), .B(n3556), .ZN(n2926) );
  XNOR2_X1 U2859 ( .A(n475), .B(n351), .ZN(n2860) );
  XNOR2_X1 U2860 ( .A(n475), .B(n363), .ZN(n2728) );
  XNOR2_X1 U2861 ( .A(n475), .B(n336), .ZN(n3025) );
  INV_X1 U2862 ( .A(n529), .ZN(n2637) );
  XNOR2_X1 U2863 ( .A(n529), .B(n366), .ZN(n2668) );
  XNOR2_X1 U2864 ( .A(n529), .B(n363), .ZN(n2701) );
  XNOR2_X1 U2865 ( .A(n529), .B(n360), .ZN(n2734) );
  XNOR2_X1 U2866 ( .A(n529), .B(n3467), .ZN(n2767) );
  XNOR2_X1 U2867 ( .A(n529), .B(n3645), .ZN(n2866) );
  XNOR2_X1 U2868 ( .A(n529), .B(n351), .ZN(n2833) );
  XNOR2_X1 U2869 ( .A(n529), .B(n354), .ZN(n2800) );
  XNOR2_X1 U2870 ( .A(n529), .B(n342), .ZN(n2932) );
  XNOR2_X1 U2871 ( .A(n529), .B(n333), .ZN(n3031) );
  XNOR2_X1 U2872 ( .A(n529), .B(n336), .ZN(n2998) );
  XNOR2_X1 U2873 ( .A(n529), .B(n339), .ZN(n2965) );
  XNOR2_X1 U2874 ( .A(n529), .B(n3502), .ZN(n3130) );
  XNOR2_X1 U2875 ( .A(n529), .B(n3556), .ZN(n2899) );
  XNOR2_X1 U2876 ( .A(n529), .B(n321), .ZN(n3163) );
  XNOR2_X1 U2877 ( .A(n529), .B(n330), .ZN(n3064) );
  XNOR2_X1 U2878 ( .A(n469), .B(n321), .ZN(n3193) );
  INV_X1 U2879 ( .A(n469), .ZN(n2667) );
  XNOR2_X1 U2880 ( .A(n469), .B(n333), .ZN(n3061) );
  XNOR2_X1 U2881 ( .A(n469), .B(n3513), .ZN(n3160) );
  XNOR2_X1 U2882 ( .A(n469), .B(n327), .ZN(n3127) );
  XNOR2_X1 U2883 ( .A(n469), .B(n336), .ZN(n3028) );
  XNOR2_X1 U2884 ( .A(n469), .B(n360), .ZN(n2764) );
  XNOR2_X1 U2885 ( .A(n469), .B(n342), .ZN(n2962) );
  XNOR2_X1 U2886 ( .A(n469), .B(n351), .ZN(n2863) );
  XNOR2_X1 U2887 ( .A(n469), .B(n354), .ZN(n2830) );
  XNOR2_X1 U2888 ( .A(n469), .B(n348), .ZN(n2896) );
  XNOR2_X1 U2889 ( .A(n469), .B(n330), .ZN(n3094) );
  XNOR2_X1 U2890 ( .A(n469), .B(n339), .ZN(n2995) );
  XNOR2_X1 U2891 ( .A(n469), .B(n366), .ZN(n2698) );
  XNOR2_X1 U2892 ( .A(n469), .B(n363), .ZN(n2731) );
  XNOR2_X1 U2893 ( .A(n469), .B(n357), .ZN(n2797) );
  XNOR2_X1 U2894 ( .A(n469), .B(n3564), .ZN(n2929) );
  XNOR2_X1 U2895 ( .A(n471), .B(n3778), .ZN(n3159) );
  XNOR2_X1 U2896 ( .A(n471), .B(n321), .ZN(n3192) );
  XNOR2_X1 U2897 ( .A(n471), .B(n333), .ZN(n3060) );
  INV_X1 U2898 ( .A(n471), .ZN(n2666) );
  XNOR2_X1 U2899 ( .A(n471), .B(n327), .ZN(n3126) );
  XNOR2_X1 U2900 ( .A(n471), .B(n330), .ZN(n3093) );
  XNOR2_X1 U2901 ( .A(n471), .B(n351), .ZN(n2862) );
  XNOR2_X1 U2902 ( .A(n471), .B(n348), .ZN(n2895) );
  XNOR2_X1 U2903 ( .A(n471), .B(n336), .ZN(n3027) );
  XNOR2_X1 U2904 ( .A(n471), .B(n342), .ZN(n2961) );
  XNOR2_X1 U2905 ( .A(n471), .B(n360), .ZN(n2763) );
  XNOR2_X1 U2906 ( .A(n471), .B(n366), .ZN(n2697) );
  XNOR2_X1 U2907 ( .A(n471), .B(n339), .ZN(n2994) );
  XNOR2_X1 U2908 ( .A(n471), .B(n354), .ZN(n2829) );
  XNOR2_X1 U2909 ( .A(n471), .B(n363), .ZN(n2730) );
  XNOR2_X1 U2910 ( .A(n471), .B(n3564), .ZN(n2928) );
  XNOR2_X1 U2911 ( .A(n471), .B(n357), .ZN(n2796) );
  INV_X1 U2912 ( .A(n527), .ZN(n2638) );
  XNOR2_X1 U2913 ( .A(n527), .B(n366), .ZN(n2669) );
  XNOR2_X1 U2914 ( .A(n527), .B(n363), .ZN(n2702) );
  XNOR2_X1 U2915 ( .A(n527), .B(n360), .ZN(n2735) );
  XNOR2_X1 U2916 ( .A(n527), .B(n3588), .ZN(n2834) );
  XNOR2_X1 U2917 ( .A(n527), .B(n357), .ZN(n2768) );
  XNOR2_X1 U2918 ( .A(n527), .B(n348), .ZN(n2867) );
  XNOR2_X1 U2919 ( .A(n527), .B(n336), .ZN(n2999) );
  XNOR2_X1 U2920 ( .A(n527), .B(n354), .ZN(n2801) );
  XNOR2_X1 U2921 ( .A(n527), .B(n3564), .ZN(n2900) );
  XNOR2_X1 U2922 ( .A(n527), .B(n327), .ZN(n3098) );
  XNOR2_X1 U2923 ( .A(n527), .B(n3502), .ZN(n3131) );
  XNOR2_X1 U2924 ( .A(n527), .B(n342), .ZN(n2933) );
  XNOR2_X1 U2925 ( .A(n527), .B(n339), .ZN(n2966) );
  XNOR2_X1 U2926 ( .A(n527), .B(n321), .ZN(n3164) );
  XNOR2_X1 U2927 ( .A(n527), .B(n330), .ZN(n3065) );
  XNOR2_X1 U2928 ( .A(n527), .B(n333), .ZN(n3032) );
  XNOR2_X1 U2929 ( .A(n473), .B(n3778), .ZN(n3158) );
  INV_X1 U2930 ( .A(n473), .ZN(n2665) );
  XNOR2_X1 U2931 ( .A(n473), .B(n333), .ZN(n3059) );
  XNOR2_X1 U2932 ( .A(n473), .B(n321), .ZN(n3191) );
  XNOR2_X1 U2933 ( .A(n473), .B(n327), .ZN(n3125) );
  XNOR2_X1 U2934 ( .A(n473), .B(n330), .ZN(n3092) );
  XNOR2_X1 U2935 ( .A(n473), .B(n351), .ZN(n2861) );
  XNOR2_X1 U2936 ( .A(n473), .B(n342), .ZN(n2960) );
  XNOR2_X1 U2937 ( .A(n473), .B(n3564), .ZN(n2927) );
  XNOR2_X1 U2938 ( .A(n473), .B(n348), .ZN(n2894) );
  XNOR2_X1 U2939 ( .A(n473), .B(n366), .ZN(n2696) );
  XNOR2_X1 U2940 ( .A(n473), .B(n360), .ZN(n2762) );
  XNOR2_X1 U2941 ( .A(n473), .B(n339), .ZN(n2993) );
  XNOR2_X1 U2942 ( .A(n473), .B(n363), .ZN(n2729) );
  XNOR2_X1 U2943 ( .A(n473), .B(n336), .ZN(n3026) );
  XNOR2_X1 U2944 ( .A(n473), .B(n354), .ZN(n2828) );
  INV_X1 U2945 ( .A(n479), .ZN(n2662) );
  XNOR2_X1 U2946 ( .A(n479), .B(n321), .ZN(n3188) );
  XNOR2_X1 U2947 ( .A(n479), .B(n3513), .ZN(n3155) );
  XNOR2_X1 U2948 ( .A(n479), .B(n354), .ZN(n2825) );
  XNOR2_X1 U2949 ( .A(n479), .B(n327), .ZN(n3122) );
  XNOR2_X1 U2950 ( .A(n479), .B(n330), .ZN(n3089) );
  XNOR2_X1 U2951 ( .A(n479), .B(n3564), .ZN(n2924) );
  XNOR2_X1 U2952 ( .A(n479), .B(n363), .ZN(n2726) );
  XNOR2_X1 U2953 ( .A(n479), .B(n336), .ZN(n3023) );
  XNOR2_X1 U2954 ( .A(n479), .B(n351), .ZN(n2858) );
  XNOR2_X1 U2955 ( .A(n479), .B(n342), .ZN(n2957) );
  XNOR2_X1 U2956 ( .A(n479), .B(n339), .ZN(n2990) );
  XNOR2_X1 U2957 ( .A(n479), .B(n348), .ZN(n2891) );
  XNOR2_X1 U2958 ( .A(n479), .B(n366), .ZN(n2693) );
  XNOR2_X1 U2959 ( .A(n479), .B(n360), .ZN(n2759) );
  XNOR2_X1 U2960 ( .A(n479), .B(n333), .ZN(n3056) );
  XNOR2_X1 U2961 ( .A(n479), .B(n357), .ZN(n2792) );
  INV_X1 U2962 ( .A(n525), .ZN(n2639) );
  XNOR2_X1 U2963 ( .A(n525), .B(n366), .ZN(n2670) );
  XNOR2_X1 U2964 ( .A(n525), .B(n363), .ZN(n2703) );
  XNOR2_X1 U2965 ( .A(n525), .B(n360), .ZN(n2736) );
  XNOR2_X1 U2966 ( .A(n525), .B(n3588), .ZN(n2835) );
  XNOR2_X1 U2967 ( .A(n525), .B(n336), .ZN(n3000) );
  XNOR2_X1 U2968 ( .A(n525), .B(n348), .ZN(n2868) );
  XNOR2_X1 U2969 ( .A(n525), .B(n354), .ZN(n2802) );
  XNOR2_X1 U2970 ( .A(n525), .B(n3564), .ZN(n2901) );
  XNOR2_X1 U2971 ( .A(n525), .B(n342), .ZN(n2934) );
  XNOR2_X1 U2972 ( .A(n525), .B(n357), .ZN(n2769) );
  XNOR2_X1 U2973 ( .A(n525), .B(n339), .ZN(n2967) );
  XNOR2_X1 U2974 ( .A(n525), .B(n3502), .ZN(n3132) );
  XNOR2_X1 U2975 ( .A(n525), .B(n330), .ZN(n3066) );
  XNOR2_X1 U2976 ( .A(n525), .B(n333), .ZN(n3033) );
  XNOR2_X1 U2977 ( .A(n525), .B(n321), .ZN(n3165) );
  INV_X1 U2978 ( .A(n523), .ZN(n2640) );
  XNOR2_X1 U2979 ( .A(n523), .B(n366), .ZN(n2671) );
  XNOR2_X1 U2980 ( .A(n523), .B(n363), .ZN(n2704) );
  XNOR2_X1 U2981 ( .A(n523), .B(n360), .ZN(n2737) );
  XNOR2_X1 U2982 ( .A(n523), .B(n354), .ZN(n2803) );
  XNOR2_X1 U2983 ( .A(n523), .B(n348), .ZN(n2869) );
  XNOR2_X1 U2984 ( .A(n523), .B(n351), .ZN(n2836) );
  XNOR2_X1 U2985 ( .A(n523), .B(n339), .ZN(n2968) );
  XNOR2_X1 U2986 ( .A(n523), .B(n357), .ZN(n2770) );
  XNOR2_X1 U2987 ( .A(n523), .B(n342), .ZN(n2935) );
  XNOR2_X1 U2988 ( .A(n523), .B(n3564), .ZN(n2902) );
  XNOR2_X1 U2989 ( .A(n523), .B(n336), .ZN(n3001) );
  XNOR2_X1 U2990 ( .A(n523), .B(n330), .ZN(n3067) );
  XNOR2_X1 U2991 ( .A(n523), .B(n3502), .ZN(n3133) );
  XNOR2_X1 U2992 ( .A(n523), .B(n333), .ZN(n3034) );
  XNOR2_X1 U2993 ( .A(n523), .B(n321), .ZN(n3166) );
  INV_X1 U2994 ( .A(n485), .ZN(n2659) );
  XNOR2_X1 U2995 ( .A(n485), .B(n321), .ZN(n3185) );
  XNOR2_X1 U2996 ( .A(n485), .B(n363), .ZN(n2723) );
  XNOR2_X1 U2997 ( .A(n485), .B(n366), .ZN(n2690) );
  XNOR2_X1 U2998 ( .A(n485), .B(n327), .ZN(n3119) );
  XNOR2_X1 U2999 ( .A(n485), .B(n3513), .ZN(n3152) );
  XNOR2_X1 U3000 ( .A(n485), .B(n354), .ZN(n2822) );
  XNOR2_X1 U3001 ( .A(n485), .B(n357), .ZN(n2789) );
  XNOR2_X1 U3002 ( .A(n485), .B(n342), .ZN(n2954) );
  XNOR2_X1 U3003 ( .A(n485), .B(n330), .ZN(n3086) );
  XNOR2_X1 U3004 ( .A(n485), .B(n351), .ZN(n2855) );
  XNOR2_X1 U3005 ( .A(n485), .B(n339), .ZN(n2987) );
  XNOR2_X1 U3006 ( .A(n485), .B(n336), .ZN(n3020) );
  XNOR2_X1 U3007 ( .A(n485), .B(n3556), .ZN(n2921) );
  XNOR2_X1 U3008 ( .A(n485), .B(n333), .ZN(n3053) );
  XNOR2_X1 U3009 ( .A(n485), .B(n360), .ZN(n2756) );
  INV_X1 U3010 ( .A(n491), .ZN(n2656) );
  XNOR2_X1 U3011 ( .A(n491), .B(n333), .ZN(n3050) );
  XNOR2_X1 U3012 ( .A(n491), .B(n363), .ZN(n2720) );
  XNOR2_X1 U3013 ( .A(n491), .B(n354), .ZN(n2819) );
  XNOR2_X1 U3014 ( .A(n491), .B(n327), .ZN(n3116) );
  XNOR2_X1 U3015 ( .A(n491), .B(n330), .ZN(n3083) );
  XNOR2_X1 U3016 ( .A(n491), .B(n366), .ZN(n2687) );
  XNOR2_X1 U3017 ( .A(n491), .B(n336), .ZN(n3017) );
  XNOR2_X1 U3018 ( .A(n491), .B(n3556), .ZN(n2918) );
  XNOR2_X1 U3019 ( .A(n491), .B(n357), .ZN(n2786) );
  XNOR2_X1 U3020 ( .A(n491), .B(n321), .ZN(n3182) );
  XNOR2_X1 U3021 ( .A(n491), .B(n342), .ZN(n2951) );
  XNOR2_X1 U3022 ( .A(n491), .B(n351), .ZN(n2852) );
  XNOR2_X1 U3023 ( .A(n491), .B(n360), .ZN(n2753) );
  XNOR2_X1 U3024 ( .A(n491), .B(n339), .ZN(n2984) );
  XNOR2_X1 U3025 ( .A(n491), .B(n324), .ZN(n3149) );
  INV_X1 U3026 ( .A(n521), .ZN(n2641) );
  XNOR2_X1 U3027 ( .A(n521), .B(n366), .ZN(n2672) );
  XNOR2_X1 U3028 ( .A(n521), .B(n363), .ZN(n2705) );
  XNOR2_X1 U3029 ( .A(n521), .B(n342), .ZN(n2936) );
  XNOR2_X1 U3030 ( .A(n521), .B(n357), .ZN(n2771) );
  XNOR2_X1 U3031 ( .A(n521), .B(n327), .ZN(n3101) );
  XNOR2_X1 U3032 ( .A(n521), .B(n354), .ZN(n2804) );
  XNOR2_X1 U3033 ( .A(n521), .B(n3564), .ZN(n2903) );
  XNOR2_X1 U3034 ( .A(n521), .B(n360), .ZN(n2738) );
  XNOR2_X1 U3035 ( .A(n521), .B(n351), .ZN(n2837) );
  XNOR2_X1 U3036 ( .A(n521), .B(n330), .ZN(n3068) );
  XNOR2_X1 U3037 ( .A(n521), .B(n348), .ZN(n2870) );
  XNOR2_X1 U3038 ( .A(n521), .B(n3502), .ZN(n3134) );
  XNOR2_X1 U3039 ( .A(n521), .B(n333), .ZN(n3035) );
  XNOR2_X1 U3040 ( .A(n521), .B(n321), .ZN(n3167) );
  XNOR2_X1 U3041 ( .A(n521), .B(n336), .ZN(n3002) );
  XNOR2_X1 U3042 ( .A(n521), .B(n339), .ZN(n2969) );
  INV_X1 U3043 ( .A(n519), .ZN(n2642) );
  XNOR2_X1 U3044 ( .A(n519), .B(n366), .ZN(n2673) );
  XNOR2_X1 U3045 ( .A(n519), .B(n363), .ZN(n2706) );
  XNOR2_X1 U3046 ( .A(n519), .B(n333), .ZN(n3036) );
  XNOR2_X1 U3047 ( .A(n519), .B(n3467), .ZN(n2772) );
  XNOR2_X1 U3048 ( .A(n519), .B(n354), .ZN(n2805) );
  XNOR2_X1 U3049 ( .A(n519), .B(n3564), .ZN(n2904) );
  XNOR2_X1 U3050 ( .A(n519), .B(n348), .ZN(n2871) );
  XNOR2_X1 U3051 ( .A(n519), .B(n360), .ZN(n2739) );
  XNOR2_X1 U3052 ( .A(n519), .B(n3634), .ZN(n2937) );
  XNOR2_X1 U3053 ( .A(n519), .B(n327), .ZN(n3102) );
  XNOR2_X1 U3054 ( .A(n519), .B(n3502), .ZN(n3135) );
  XNOR2_X1 U3055 ( .A(n519), .B(n351), .ZN(n2838) );
  XNOR2_X1 U3056 ( .A(n519), .B(n330), .ZN(n3069) );
  XNOR2_X1 U3057 ( .A(n519), .B(n336), .ZN(n3003) );
  XNOR2_X1 U3058 ( .A(n519), .B(n321), .ZN(n3168) );
  XNOR2_X1 U3059 ( .A(n519), .B(n339), .ZN(n2970) );
  INV_X1 U3060 ( .A(n517), .ZN(n2643) );
  XNOR2_X1 U3061 ( .A(n517), .B(n366), .ZN(n2674) );
  XNOR2_X1 U3062 ( .A(n517), .B(n363), .ZN(n2707) );
  XNOR2_X1 U3063 ( .A(n517), .B(n3467), .ZN(n2773) );
  XNOR2_X1 U3064 ( .A(n517), .B(n333), .ZN(n3037) );
  XNOR2_X1 U3065 ( .A(n517), .B(n360), .ZN(n2740) );
  XNOR2_X1 U3066 ( .A(n517), .B(n3564), .ZN(n2905) );
  XNOR2_X1 U3067 ( .A(n517), .B(n348), .ZN(n2872) );
  XNOR2_X1 U3068 ( .A(n517), .B(n351), .ZN(n2839) );
  XNOR2_X1 U3069 ( .A(n517), .B(n327), .ZN(n3103) );
  XNOR2_X1 U3070 ( .A(n517), .B(n3502), .ZN(n3136) );
  XNOR2_X1 U3071 ( .A(n517), .B(n354), .ZN(n2806) );
  XNOR2_X1 U3072 ( .A(n517), .B(n336), .ZN(n3004) );
  XNOR2_X1 U3073 ( .A(n517), .B(n330), .ZN(n3070) );
  XNOR2_X1 U3074 ( .A(n517), .B(n342), .ZN(n2938) );
  XNOR2_X1 U3075 ( .A(n517), .B(n339), .ZN(n2971) );
  XNOR2_X1 U3076 ( .A(n517), .B(n321), .ZN(n3169) );
  INV_X1 U3077 ( .A(n497), .ZN(n2653) );
  XNOR2_X1 U3078 ( .A(n497), .B(n366), .ZN(n2684) );
  XNOR2_X1 U3079 ( .A(n497), .B(n357), .ZN(n2783) );
  XNOR2_X1 U3080 ( .A(n497), .B(n360), .ZN(n2750) );
  XNOR2_X1 U3081 ( .A(n497), .B(n348), .ZN(n2882) );
  XNOR2_X1 U3082 ( .A(n497), .B(n333), .ZN(n3047) );
  XNOR2_X1 U3083 ( .A(n497), .B(n363), .ZN(n2717) );
  XNOR2_X1 U3084 ( .A(n497), .B(n327), .ZN(n3113) );
  XNOR2_X1 U3085 ( .A(n497), .B(n3502), .ZN(n3146) );
  XNOR2_X1 U3086 ( .A(n497), .B(n342), .ZN(n2948) );
  XNOR2_X1 U3087 ( .A(n497), .B(n351), .ZN(n2849) );
  XNOR2_X1 U3088 ( .A(n497), .B(n3556), .ZN(n2915) );
  XNOR2_X1 U3089 ( .A(n497), .B(n330), .ZN(n3080) );
  XNOR2_X1 U3090 ( .A(n497), .B(n336), .ZN(n3014) );
  XNOR2_X1 U3091 ( .A(n497), .B(n339), .ZN(n2981) );
  XNOR2_X1 U3092 ( .A(n497), .B(n354), .ZN(n2816) );
  XNOR2_X1 U3093 ( .A(n497), .B(n321), .ZN(n3179) );
  INV_X1 U3094 ( .A(n503), .ZN(n2650) );
  XNOR2_X1 U3095 ( .A(n503), .B(n327), .ZN(n3110) );
  XNOR2_X1 U3096 ( .A(n503), .B(n366), .ZN(n2681) );
  XNOR2_X1 U3097 ( .A(n503), .B(n342), .ZN(n2945) );
  XNOR2_X1 U3098 ( .A(n503), .B(n363), .ZN(n2714) );
  XNOR2_X1 U3099 ( .A(n503), .B(n354), .ZN(n2813) );
  XNOR2_X1 U3100 ( .A(n503), .B(n357), .ZN(n2780) );
  XNOR2_X1 U3101 ( .A(n503), .B(n351), .ZN(n2846) );
  XNOR2_X1 U3102 ( .A(n503), .B(n3556), .ZN(n2912) );
  XNOR2_X1 U3103 ( .A(n503), .B(n339), .ZN(n2978) );
  XNOR2_X1 U3104 ( .A(n503), .B(n360), .ZN(n2747) );
  XNOR2_X1 U3105 ( .A(n503), .B(n333), .ZN(n3044) );
  XNOR2_X1 U3106 ( .A(n503), .B(n324), .ZN(n3143) );
  XNOR2_X1 U3107 ( .A(n503), .B(n330), .ZN(n3077) );
  XNOR2_X1 U3108 ( .A(n503), .B(n336), .ZN(n3011) );
  XNOR2_X1 U3109 ( .A(n503), .B(n348), .ZN(n2879) );
  XNOR2_X1 U3110 ( .A(n503), .B(n321), .ZN(n3176) );
  INV_X1 U3111 ( .A(n515), .ZN(n2644) );
  XNOR2_X1 U3112 ( .A(n515), .B(n363), .ZN(n2708) );
  XNOR2_X1 U3113 ( .A(n515), .B(n366), .ZN(n2675) );
  XNOR2_X1 U3114 ( .A(n515), .B(n3467), .ZN(n2774) );
  XNOR2_X1 U3115 ( .A(n515), .B(n360), .ZN(n2741) );
  XNOR2_X1 U3116 ( .A(n515), .B(n3564), .ZN(n2906) );
  XNOR2_X1 U3117 ( .A(n515), .B(n351), .ZN(n2840) );
  XNOR2_X1 U3118 ( .A(n515), .B(n327), .ZN(n3104) );
  XNOR2_X1 U3119 ( .A(n515), .B(n354), .ZN(n2807) );
  XNOR2_X1 U3120 ( .A(n515), .B(n348), .ZN(n2873) );
  XNOR2_X1 U3121 ( .A(n515), .B(n336), .ZN(n3005) );
  XNOR2_X1 U3122 ( .A(n515), .B(n330), .ZN(n3071) );
  XNOR2_X1 U3123 ( .A(n515), .B(n3502), .ZN(n3137) );
  XNOR2_X1 U3124 ( .A(n515), .B(n342), .ZN(n2939) );
  XNOR2_X1 U3125 ( .A(n515), .B(n333), .ZN(n3038) );
  XNOR2_X1 U3126 ( .A(n515), .B(n339), .ZN(n2972) );
  XNOR2_X1 U3127 ( .A(n515), .B(n321), .ZN(n3170) );
  INV_X1 U3128 ( .A(n509), .ZN(n2647) );
  XNOR2_X1 U3129 ( .A(n509), .B(n363), .ZN(n2711) );
  XNOR2_X1 U3130 ( .A(n509), .B(n330), .ZN(n3074) );
  XNOR2_X1 U3131 ( .A(n509), .B(n366), .ZN(n2678) );
  XNOR2_X1 U3132 ( .A(n509), .B(n357), .ZN(n2777) );
  XNOR2_X1 U3133 ( .A(n509), .B(n360), .ZN(n2744) );
  XNOR2_X1 U3134 ( .A(n509), .B(n351), .ZN(n2843) );
  XNOR2_X1 U3135 ( .A(n509), .B(n3502), .ZN(n3140) );
  XNOR2_X1 U3136 ( .A(n509), .B(n342), .ZN(n2942) );
  XNOR2_X1 U3137 ( .A(n509), .B(n354), .ZN(n2810) );
  XNOR2_X1 U3138 ( .A(n509), .B(n333), .ZN(n3041) );
  XNOR2_X1 U3139 ( .A(n509), .B(n336), .ZN(n3008) );
  XNOR2_X1 U3140 ( .A(n509), .B(n321), .ZN(n3173) );
  XNOR2_X1 U3141 ( .A(n509), .B(n339), .ZN(n2975) );
  XNOR2_X1 U3142 ( .A(n509), .B(n345), .ZN(n2909) );
  NAND2_X1 U3143 ( .A1(n851), .A2(n850), .ZN(n571) );
  OAI21_X1 U3144 ( .B1(n855), .B2(n849), .A(n850), .ZN(n848) );
  NAND2_X1 U3145 ( .A1(n1798), .A2(n1819), .ZN(n850) );
  NOR2_X1 U3146 ( .A1(n1798), .A2(n1819), .ZN(n849) );
  INV_X2 U3147 ( .A(a[6]), .ZN(n3701) );
  INV_X2 U3148 ( .A(n3647), .ZN(n3648) );
  INV_X2 U3149 ( .A(n3647), .ZN(n3650) );
  NOR2_X2 U3150 ( .A1(n1750), .A2(n1773), .ZN(n839) );
  INV_X1 U3151 ( .A(n3416), .ZN(n3635) );
  AOI21_X1 U3152 ( .B1(n832), .B2(n838), .A(n833), .ZN(n3409) );
  AOI21_X1 U3153 ( .B1(n832), .B2(n838), .A(n833), .ZN(n831) );
  INV_X2 U3154 ( .A(n3636), .ZN(n3638) );
  INV_X2 U3155 ( .A(n3636), .ZN(n3639) );
  INV_X1 U3156 ( .A(n3521), .ZN(n3636) );
  INV_X1 U3157 ( .A(n846), .ZN(n844) );
  XOR2_X1 U3158 ( .A(n1821), .B(n1802), .Z(n3410) );
  XOR2_X1 U3159 ( .A(n1800), .B(n3410), .Z(n1798) );
  NAND2_X1 U3160 ( .A1(n1800), .A2(n1821), .ZN(n3411) );
  NAND2_X1 U3161 ( .A1(n1800), .A2(n1802), .ZN(n3412) );
  NAND2_X1 U3162 ( .A1(n1821), .A2(n1802), .ZN(n3413) );
  NAND3_X1 U3163 ( .A1(n3411), .A2(n3413), .A3(n3412), .ZN(n1797) );
  AOI21_X1 U3164 ( .B1(n749), .B2(n999), .A(n746), .ZN(n3414) );
  AOI21_X1 U3165 ( .B1(n749), .B2(n999), .A(n746), .ZN(n744) );
  BUF_X1 U3166 ( .A(n612), .Z(n3415) );
  AOI21_X2 U3167 ( .B1(n612), .B2(n981), .A(n607), .ZN(n605) );
  OAI21_X2 U3168 ( .B1(n777), .B2(n781), .A(n778), .ZN(n776) );
  XNOR2_X1 U3169 ( .A(n3489), .B(n327), .ZN(n3241) );
  INV_X4 U3170 ( .A(a[4]), .ZN(n3489) );
  AOI21_X1 U3171 ( .B1(n878), .B2(n897), .A(n879), .ZN(n877) );
  OAI21_X2 U3172 ( .B1(n898), .B2(n915), .A(n899), .ZN(n897) );
  NAND2_X1 U3173 ( .A1(n905), .A2(n900), .ZN(n898) );
  AOI21_X2 U3174 ( .B1(n906), .B2(n900), .A(n901), .ZN(n899) );
  OAI22_X1 U3175 ( .A1(n3551), .A2(n2808), .B1(n2807), .B2(n3469), .ZN(n2239)
         );
  OAI22_X1 U3176 ( .A1(n3551), .A2(n2813), .B1(n2812), .B2(n3469), .ZN(n2244)
         );
  OAI22_X1 U3177 ( .A1(n3551), .A2(n2809), .B1(n2808), .B2(n3469), .ZN(n2240)
         );
  OAI22_X1 U3178 ( .A1(n3551), .A2(n2803), .B1(n2802), .B2(n3469), .ZN(n2234)
         );
  OAI22_X1 U3179 ( .A1(n3551), .A2(n2800), .B1(n3469), .B2(n3281), .ZN(n2231)
         );
  OAI22_X1 U3180 ( .A1(n3551), .A2(n2824), .B1(n2823), .B2(n3469), .ZN(n2255)
         );
  OAI22_X1 U3181 ( .A1(n3551), .A2(n2831), .B1(n2830), .B2(n3469), .ZN(n2262)
         );
  OAI22_X1 U3182 ( .A1(n3551), .A2(n2825), .B1(n2824), .B2(n3469), .ZN(n2256)
         );
  OAI22_X1 U3183 ( .A1(n3551), .A2(n2826), .B1(n2825), .B2(n3469), .ZN(n2257)
         );
  OAI22_X1 U3184 ( .A1(n3551), .A2(n2828), .B1(n2827), .B2(n3469), .ZN(n2259)
         );
  OAI22_X1 U3185 ( .A1(n3551), .A2(n2811), .B1(n2810), .B2(n3469), .ZN(n2242)
         );
  OAI22_X1 U3186 ( .A1(n3551), .A2(n2810), .B1(n2809), .B2(n3469), .ZN(n2241)
         );
  OR2_X4 U3187 ( .A1(n3417), .A2(n3757), .ZN(n3416) );
  XOR2_X2 U3188 ( .A(n3457), .B(n339), .Z(n3417) );
  OAI21_X1 U3189 ( .B1(n819), .B2(n825), .A(n820), .ZN(n3418) );
  OAI21_X1 U3190 ( .B1(n819), .B2(n825), .A(n820), .ZN(n818) );
  AOI21_X1 U3191 ( .B1(n885), .B2(n893), .A(n886), .ZN(n3419) );
  AOI21_X1 U3192 ( .B1(n885), .B2(n893), .A(n886), .ZN(n884) );
  INV_X1 U3193 ( .A(n1005), .ZN(n3420) );
  INV_X2 U3194 ( .A(n3671), .ZN(n3456) );
  OAI22_X1 U3195 ( .A1(n3552), .A2(n2816), .B1(n2815), .B2(n3469), .ZN(n2247)
         );
  OAI22_X1 U3196 ( .A1(n3552), .A2(n2820), .B1(n2819), .B2(n3469), .ZN(n2251)
         );
  OAI22_X1 U3197 ( .A1(n3552), .A2(n2804), .B1(n2803), .B2(n3469), .ZN(n2235)
         );
  OAI22_X1 U3198 ( .A1(n3552), .A2(n2814), .B1(n2813), .B2(n3469), .ZN(n2245)
         );
  OAI22_X1 U3199 ( .A1(n3552), .A2(n3281), .B1(n2832), .B2(n3469), .ZN(n2065)
         );
  OAI22_X1 U3200 ( .A1(n3552), .A2(n2801), .B1(n2800), .B2(n3469), .ZN(n2232)
         );
  OAI22_X1 U3201 ( .A1(n3552), .A2(n2806), .B1(n2805), .B2(n3469), .ZN(n2237)
         );
  OAI22_X1 U3202 ( .A1(n3552), .A2(n2802), .B1(n2801), .B2(n3469), .ZN(n2233)
         );
  OAI22_X1 U3203 ( .A1(n3552), .A2(n2812), .B1(n2811), .B2(n3469), .ZN(n2243)
         );
  OAI22_X1 U3204 ( .A1(n3552), .A2(n2827), .B1(n2826), .B2(n3469), .ZN(n2258)
         );
  OAI22_X1 U3205 ( .A1(n3552), .A2(n2807), .B1(n2806), .B2(n3469), .ZN(n2238)
         );
  OAI22_X1 U3206 ( .A1(n3552), .A2(n2805), .B1(n2804), .B2(n3469), .ZN(n2236)
         );
  OAI22_X1 U3207 ( .A1(n3552), .A2(n2829), .B1(n2828), .B2(n3469), .ZN(n2260)
         );
  INV_X1 U3208 ( .A(n888), .ZN(n886) );
  OAI21_X1 U3209 ( .B1(n855), .B2(n842), .A(n843), .ZN(n841) );
  OAI22_X1 U3210 ( .A1(n3416), .A2(n2982), .B1(n2981), .B2(n387), .ZN(n2418)
         );
  XNOR2_X1 U3211 ( .A(n3421), .B(n1535), .ZN(n1527) );
  XNOR2_X1 U3212 ( .A(n1562), .B(n1537), .ZN(n3421) );
  NAND2_X1 U3213 ( .A1(n3422), .A2(n3423), .ZN(n3424) );
  NAND2_X1 U3214 ( .A1(n3424), .A2(n858), .ZN(n856) );
  INV_X1 U3215 ( .A(n877), .ZN(n3422) );
  INV_X1 U3216 ( .A(n857), .ZN(n3423) );
  BUF_X1 U3217 ( .A(a[18]), .Z(n3425) );
  XOR2_X2 U3218 ( .A(n1584), .B(n3515), .Z(n1582) );
  INV_X2 U3219 ( .A(n3688), .ZN(n440) );
  XNOR2_X2 U3220 ( .A(n3752), .B(n3288), .ZN(n3426) );
  INV_X4 U3221 ( .A(n3426), .ZN(n3751) );
  INV_X4 U3222 ( .A(n333), .ZN(n3288) );
  NAND2_X2 U3223 ( .A1(n3455), .A2(n360), .ZN(n3616) );
  NAND2_X2 U3224 ( .A1(n1519), .A2(n1550), .ZN(n794) );
  XOR2_X1 U3225 ( .A(n3755), .B(n3279), .Z(n3230) );
  INV_X4 U3226 ( .A(n360), .ZN(n3279) );
  BUF_X1 U3227 ( .A(n815), .Z(n3427) );
  INV_X2 U3228 ( .A(n3688), .ZN(n3580) );
  XOR2_X1 U3229 ( .A(n1721), .B(n1715), .Z(n3428) );
  XOR2_X1 U3230 ( .A(n3428), .B(n1719), .Z(n1684) );
  XOR2_X1 U3231 ( .A(n1707), .B(n1682), .Z(n3429) );
  XOR2_X1 U3232 ( .A(n3429), .B(n1684), .Z(n1676) );
  NAND2_X1 U3233 ( .A1(n1721), .A2(n1715), .ZN(n3430) );
  NAND2_X1 U3234 ( .A1(n1721), .A2(n1719), .ZN(n3431) );
  NAND2_X1 U3235 ( .A1(n1715), .A2(n1719), .ZN(n3432) );
  NAND3_X1 U3236 ( .A1(n3430), .A2(n3431), .A3(n3432), .ZN(n1683) );
  NAND2_X1 U3237 ( .A1(n1707), .A2(n1682), .ZN(n3433) );
  NAND2_X1 U3238 ( .A1(n1707), .A2(n1684), .ZN(n3434) );
  NAND2_X1 U3239 ( .A1(n1682), .A2(n1684), .ZN(n3435) );
  NAND3_X1 U3240 ( .A1(n3433), .A2(n3434), .A3(n3435), .ZN(n1675) );
  OR2_X1 U3241 ( .A1(n3562), .A2(n2888), .ZN(n3436) );
  OR2_X1 U3242 ( .A1(n2887), .A2(n396), .ZN(n3437) );
  NAND2_X1 U3243 ( .A1(n3436), .A2(n3437), .ZN(n2321) );
  XNOR2_X1 U3244 ( .A(n485), .B(n348), .ZN(n2888) );
  XNOR2_X1 U3245 ( .A(n487), .B(n348), .ZN(n2887) );
  AND2_X1 U3246 ( .A1(n3232), .A2(n3469), .ZN(n3661) );
  NAND2_X1 U3247 ( .A1(n994), .A2(n705), .ZN(n548) );
  NAND2_X1 U3248 ( .A1(n690), .A2(n615), .ZN(n613) );
  INV_X1 U3249 ( .A(n690), .ZN(n688) );
  NAND2_X1 U3250 ( .A1(n694), .A2(n994), .ZN(n692) );
  BUF_X1 U3251 ( .A(n3290), .Z(n3438) );
  NOR2_X2 U3252 ( .A1(n780), .A2(n777), .ZN(n775) );
  XNOR2_X1 U3253 ( .A(n1433), .B(n3439), .ZN(n1431) );
  XNOR2_X1 U3254 ( .A(n1460), .B(n1435), .ZN(n3439) );
  XOR2_X1 U3255 ( .A(n1409), .B(n1436), .Z(n3440) );
  XOR2_X1 U3256 ( .A(n1434), .B(n3440), .Z(n1405) );
  NAND2_X1 U3257 ( .A1(n1434), .A2(n1409), .ZN(n3441) );
  NAND2_X1 U3258 ( .A1(n1434), .A2(n1436), .ZN(n3442) );
  NAND2_X1 U3259 ( .A1(n1409), .A2(n1436), .ZN(n3443) );
  NAND3_X1 U3260 ( .A1(n3441), .A2(n3443), .A3(n3442), .ZN(n1404) );
  OAI22_X1 U3261 ( .A1(n3561), .A2(n2879), .B1(n2878), .B2(n396), .ZN(n2312)
         );
  AOI21_X1 U3262 ( .B1(n726), .B2(n709), .A(n710), .ZN(n708) );
  INV_X1 U3263 ( .A(n760), .ZN(n758) );
  AOI21_X1 U3264 ( .B1(n635), .B2(n676), .A(n636), .ZN(n634) );
  OAI21_X1 U3265 ( .B1(n634), .B2(n617), .A(n618), .ZN(n616) );
  INV_X1 U3266 ( .A(n634), .ZN(n632) );
  INV_X2 U3267 ( .A(n3763), .ZN(n428) );
  OAI21_X1 U3268 ( .B1(n3503), .B2(n857), .A(n858), .ZN(n3690) );
  XNOR2_X1 U3269 ( .A(n3752), .B(n336), .ZN(n3544) );
  XNOR2_X1 U3270 ( .A(n1405), .B(n3444), .ZN(n1403) );
  XNOR2_X1 U3271 ( .A(n1432), .B(n1407), .ZN(n3444) );
  INV_X2 U3272 ( .A(n3761), .ZN(n390) );
  XOR2_X1 U3273 ( .A(n1364), .B(n1347), .Z(n3445) );
  XOR2_X1 U3274 ( .A(n3445), .B(n1362), .Z(n1335) );
  XOR2_X1 U3275 ( .A(n1358), .B(n1337), .Z(n3446) );
  XOR2_X1 U3276 ( .A(n3446), .B(n1335), .Z(n1331) );
  NAND2_X1 U3277 ( .A1(n1364), .A2(n1347), .ZN(n3447) );
  NAND2_X1 U3278 ( .A1(n1364), .A2(n1362), .ZN(n3448) );
  NAND2_X1 U3279 ( .A1(n1347), .A2(n1362), .ZN(n3449) );
  NAND3_X1 U3280 ( .A1(n3447), .A2(n3448), .A3(n3449), .ZN(n1334) );
  NAND2_X1 U3281 ( .A1(n1358), .A2(n1337), .ZN(n3450) );
  NAND2_X1 U3282 ( .A1(n1358), .A2(n1335), .ZN(n3451) );
  NAND2_X1 U3283 ( .A1(n1337), .A2(n1335), .ZN(n3452) );
  NAND3_X1 U3284 ( .A1(n3450), .A2(n3451), .A3(n3452), .ZN(n1330) );
  OR2_X1 U3285 ( .A1(n446), .A2(n2877), .ZN(n3453) );
  OR2_X1 U3286 ( .A1(n2876), .A2(n396), .ZN(n3454) );
  NAND2_X1 U3287 ( .A1(n3453), .A2(n3454), .ZN(n2310) );
  XNOR2_X1 U3288 ( .A(n507), .B(n348), .ZN(n2877) );
  XNOR2_X1 U3289 ( .A(n509), .B(n348), .ZN(n2876) );
  OAI22_X1 U3290 ( .A1(n440), .A2(n2944), .B1(n2943), .B2(n3649), .ZN(n2379)
         );
  OAI22_X1 U3291 ( .A1(n440), .A2(n2937), .B1(n2936), .B2(n3649), .ZN(n2372)
         );
  OAI22_X1 U3292 ( .A1(n440), .A2(n2955), .B1(n2954), .B2(n3650), .ZN(n2390)
         );
  OAI22_X1 U3293 ( .A1(n440), .A2(n3285), .B1(n2964), .B2(n3650), .ZN(n2069)
         );
  OAI22_X1 U3294 ( .A1(n3579), .A2(n2938), .B1(n2937), .B2(n3650), .ZN(n2373)
         );
  OAI22_X1 U3295 ( .A1(n3579), .A2(n2958), .B1(n2957), .B2(n3650), .ZN(n2393)
         );
  OAI22_X1 U3296 ( .A1(n440), .A2(n2933), .B1(n2932), .B2(n3649), .ZN(n2368)
         );
  OAI22_X1 U3297 ( .A1(n3579), .A2(n2945), .B1(n2944), .B2(n3650), .ZN(n2380)
         );
  OAI22_X1 U3298 ( .A1(n3579), .A2(n2960), .B1(n2959), .B2(n3649), .ZN(n2395)
         );
  OAI22_X1 U3299 ( .A1(n440), .A2(n2948), .B1(n2947), .B2(n3649), .ZN(n2383)
         );
  OAI22_X1 U3300 ( .A1(n3579), .A2(n2941), .B1(n2940), .B2(n3650), .ZN(n2376)
         );
  OAI22_X1 U3301 ( .A1(n3579), .A2(n2962), .B1(n2961), .B2(n3650), .ZN(n2397)
         );
  OAI22_X1 U3302 ( .A1(n3579), .A2(n2940), .B1(n2939), .B2(n3650), .ZN(n2375)
         );
  OAI22_X1 U3303 ( .A1(n3579), .A2(n2951), .B1(n2950), .B2(n3650), .ZN(n2386)
         );
  OAI22_X1 U3304 ( .A1(n3579), .A2(n2932), .B1(n3650), .B2(n3285), .ZN(n2367)
         );
  NOR2_X2 U3305 ( .A1(n1259), .A2(n1280), .ZN(n735) );
  AND2_X2 U3306 ( .A1(n3544), .A2(n3426), .ZN(n3543) );
  INV_X1 U3307 ( .A(n819), .ZN(n1012) );
  INV_X4 U3308 ( .A(a[28]), .ZN(n3455) );
  INV_X2 U3309 ( .A(a[28]), .ZN(n3754) );
  OAI22_X1 U3310 ( .A1(n428), .A2(n3067), .B1(n3066), .B2(n3604), .ZN(n2506)
         );
  XNOR2_X2 U3311 ( .A(n3762), .B(n339), .ZN(n3761) );
  INV_X4 U3312 ( .A(n3688), .ZN(n3579) );
  OAI22_X1 U3313 ( .A1(n3580), .A2(n2942), .B1(n2941), .B2(n3650), .ZN(n2377)
         );
  NOR2_X1 U3314 ( .A1(n3630), .A2(n613), .ZN(n611) );
  XNOR2_X2 U3315 ( .A(n3509), .B(n1521), .ZN(n1519) );
  INV_X4 U3316 ( .A(a[12]), .ZN(n3457) );
  AND2_X2 U3317 ( .A1(n3234), .A2(n396), .ZN(n3764) );
  BUF_X1 U3318 ( .A(n738), .Z(n3458) );
  AND2_X4 U3319 ( .A1(n3240), .A2(n3603), .ZN(n3763) );
  INV_X2 U3320 ( .A(n455), .ZN(n3459) );
  INV_X1 U3321 ( .A(n3459), .ZN(n3460) );
  INV_X4 U3322 ( .A(n3459), .ZN(n3462) );
  INV_X4 U3323 ( .A(n3459), .ZN(n3461) );
  INV_X1 U3324 ( .A(n735), .ZN(n997) );
  NAND2_X1 U3325 ( .A1(n998), .A2(n997), .ZN(n731) );
  OAI21_X1 U3326 ( .B1(n692), .B2(n712), .A(n693), .ZN(n691) );
  NOR2_X1 U3327 ( .A1(n1219), .A2(n1238), .ZN(n715) );
  NAND2_X1 U3328 ( .A1(n1219), .A2(n1238), .ZN(n716) );
  INV_X1 U3329 ( .A(n3671), .ZN(n3660) );
  XOR2_X1 U3330 ( .A(n3481), .B(n366), .Z(n3228) );
  NOR2_X1 U3331 ( .A1(n1377), .A2(n1402), .ZN(n3463) );
  FA_X1 U3332 ( .A(n1404), .B(n1381), .CI(n1379), .S(n3464) );
  NOR2_X1 U3333 ( .A1(n1377), .A2(n1402), .ZN(n769) );
  BUF_X1 U3334 ( .A(n781), .Z(n3465) );
  INV_X2 U3335 ( .A(n357), .ZN(n3466) );
  INV_X1 U3336 ( .A(n3467), .ZN(n3280) );
  AND2_X1 U3337 ( .A1(n3586), .A2(n3587), .ZN(n3468) );
  AND2_X4 U3338 ( .A1(n3586), .A2(n3587), .ZN(n3469) );
  BUF_X1 U3339 ( .A(n753), .Z(n3470) );
  XNOR2_X1 U3340 ( .A(a[24]), .B(n357), .ZN(n3589) );
  NAND2_X4 U3341 ( .A1(n3677), .A2(n3678), .ZN(n3704) );
  NAND2_X4 U3342 ( .A1(n3682), .A2(n3683), .ZN(n3699) );
  NAND2_X2 U3343 ( .A1(a[18]), .A2(n3681), .ZN(n3682) );
  INV_X1 U3344 ( .A(n3649), .ZN(n3471) );
  INV_X4 U3345 ( .A(n3647), .ZN(n3649) );
  AND2_X2 U3346 ( .A1(n3242), .A2(n3601), .ZN(n3672) );
  NAND2_X1 U3347 ( .A1(n611), .A2(n981), .ZN(n604) );
  NAND2_X1 U3348 ( .A1(n1005), .A2(n3465), .ZN(n559) );
  NAND2_X1 U3349 ( .A1(n1459), .A2(n1488), .ZN(n781) );
  XOR2_X1 U3350 ( .A(n2385), .B(n2449), .Z(n3472) );
  XOR2_X2 U3351 ( .A(n3472), .B(n2417), .Z(n1714) );
  XOR2_X1 U3352 ( .A(n1741), .B(n1739), .Z(n3473) );
  XOR2_X1 U3353 ( .A(n3473), .B(n1714), .Z(n1710) );
  NAND2_X1 U3354 ( .A1(n3480), .A2(n2449), .ZN(n3474) );
  NAND2_X1 U3355 ( .A1(n3480), .A2(n2417), .ZN(n3475) );
  NAND2_X2 U3356 ( .A1(n2449), .A2(n2417), .ZN(n3476) );
  NAND3_X1 U3357 ( .A1(n3474), .A2(n3475), .A3(n3476), .ZN(n1713) );
  NAND2_X1 U3358 ( .A1(n1741), .A2(n1739), .ZN(n3477) );
  NAND2_X1 U3359 ( .A1(n1741), .A2(n1714), .ZN(n3478) );
  NAND2_X1 U3360 ( .A1(n1739), .A2(n1714), .ZN(n3479) );
  NAND3_X1 U3361 ( .A1(n3477), .A2(n3478), .A3(n3479), .ZN(n1709) );
  BUF_X1 U3362 ( .A(n2385), .Z(n3480) );
  NAND2_X1 U3363 ( .A1(n3739), .A2(n363), .ZN(n3483) );
  NAND2_X1 U3364 ( .A1(n3481), .A2(n3482), .ZN(n3484) );
  NAND2_X1 U3365 ( .A1(n3483), .A2(n3484), .ZN(n3738) );
  INV_X1 U3366 ( .A(n3739), .ZN(n3481) );
  NAND2_X1 U3367 ( .A1(n1000), .A2(n755), .ZN(n554) );
  NAND2_X2 U3368 ( .A1(n3629), .A2(n351), .ZN(n3586) );
  AND2_X2 U3369 ( .A1(n3229), .A2(n411), .ZN(n3671) );
  INV_X4 U3370 ( .A(n3671), .ZN(n461) );
  NAND2_X4 U3371 ( .A1(n3680), .A2(n345), .ZN(n3683) );
  NOR2_X1 U3372 ( .A1(n784), .A2(n765), .ZN(n3486) );
  NOR2_X1 U3373 ( .A1(n784), .A2(n765), .ZN(n3485) );
  NAND2_X2 U3374 ( .A1(n3520), .A2(n775), .ZN(n765) );
  INV_X1 U3375 ( .A(n375), .ZN(n3487) );
  INV_X4 U3376 ( .A(n3487), .ZN(n3488) );
  INV_X1 U3377 ( .A(n3489), .ZN(n3490) );
  NOR2_X2 U3378 ( .A1(n3630), .A2(n688), .ZN(n686) );
  NOR2_X1 U3379 ( .A1(n788), .A2(n793), .ZN(n3491) );
  NOR2_X1 U3380 ( .A1(n788), .A2(n793), .ZN(n786) );
  NAND2_X1 U3381 ( .A1(n1405), .A2(n1432), .ZN(n3492) );
  NAND2_X1 U3382 ( .A1(n1405), .A2(n1407), .ZN(n3493) );
  NAND2_X1 U3383 ( .A1(n1432), .A2(n1407), .ZN(n3494) );
  NAND3_X1 U3384 ( .A1(n3492), .A2(n3494), .A3(n3493), .ZN(n1402) );
  NOR2_X2 U3385 ( .A1(n1724), .A2(n1749), .ZN(n834) );
  NOR2_X2 U3386 ( .A1(n3495), .A2(n3766), .ZN(n3679) );
  XNOR2_X1 U3387 ( .A(a[8]), .B(n333), .ZN(n3495) );
  OAI21_X1 U3388 ( .B1(n3606), .B2(n794), .A(n789), .ZN(n787) );
  OAI22_X1 U3389 ( .A1(n3653), .A2(n2669), .B1(n2668), .B2(n3626), .ZN(n2096)
         );
  OAI22_X1 U3390 ( .A1(n3653), .A2(n2672), .B1(n2671), .B2(n3626), .ZN(n2099)
         );
  OAI22_X1 U3391 ( .A1(n3653), .A2(n2674), .B1(n2673), .B2(n3626), .ZN(n2101)
         );
  NOR2_X1 U3392 ( .A1(n3626), .A2(n3784), .ZN(n2127) );
  OAI21_X1 U3393 ( .B1(n728), .B2(n688), .A(n689), .ZN(n3496) );
  BUF_X1 U3394 ( .A(n754), .Z(n3497) );
  OAI21_X1 U3395 ( .B1(n728), .B2(n688), .A(n689), .ZN(n687) );
  BUF_X1 U3396 ( .A(n425), .Z(n3498) );
  INV_X2 U3397 ( .A(n416), .ZN(n3499) );
  INV_X16 U3398 ( .A(n3499), .ZN(n3500) );
  OAI22_X1 U3399 ( .A1(n3416), .A2(n2976), .B1(n2975), .B2(n387), .ZN(n2412)
         );
  AOI21_X1 U3400 ( .B1(n878), .B2(n897), .A(n3506), .ZN(n3504) );
  AOI21_X1 U3401 ( .B1(n878), .B2(n897), .A(n3505), .ZN(n3503) );
  OAI21_X1 U3402 ( .B1(n3419), .B2(n880), .A(n881), .ZN(n3506) );
  OAI21_X1 U3403 ( .B1(n3419), .B2(n880), .A(n881), .ZN(n3505) );
  BUF_X1 U3404 ( .A(n425), .Z(n3507) );
  OAI21_X1 U3405 ( .B1(n884), .B2(n880), .A(n881), .ZN(n879) );
  AOI21_X2 U3406 ( .B1(n3690), .B2(n828), .A(n3720), .ZN(n3719) );
  AOI21_X1 U3407 ( .B1(n603), .B2(n980), .A(n600), .ZN(n3508) );
  AOI21_X1 U3408 ( .B1(n603), .B2(n980), .A(n600), .ZN(n598) );
  XOR2_X1 U3409 ( .A(n774), .B(n557), .Z(product[38]) );
  OAI21_X1 U3410 ( .B1(n701), .B2(n699), .A(n700), .ZN(n698) );
  XNOR2_X1 U3411 ( .A(n1552), .B(n1523), .ZN(n3509) );
  INV_X1 U3412 ( .A(n3470), .ZN(n751) );
  INV_X1 U3413 ( .A(n3759), .ZN(n3510) );
  XOR2_X1 U3414 ( .A(a[20]), .B(n351), .Z(n3233) );
  OAI22_X1 U3415 ( .A1(n3562), .A2(n2867), .B1(n2866), .B2(n396), .ZN(n2300)
         );
  OAI22_X1 U3416 ( .A1(n3562), .A2(n2876), .B1(n2875), .B2(n396), .ZN(n2309)
         );
  OAI22_X1 U3417 ( .A1(n3561), .A2(n2883), .B1(n2882), .B2(n396), .ZN(n2316)
         );
  OAI22_X1 U3418 ( .A1(n3562), .A2(n2873), .B1(n2872), .B2(n396), .ZN(n2306)
         );
  OAI22_X1 U3419 ( .A1(n3561), .A2(n2892), .B1(n2891), .B2(n396), .ZN(n2325)
         );
  OAI22_X1 U3420 ( .A1(n3562), .A2(n2874), .B1(n2873), .B2(n396), .ZN(n2307)
         );
  OAI22_X1 U3421 ( .A1(n3561), .A2(n2889), .B1(n2888), .B2(n396), .ZN(n2322)
         );
  OAI22_X1 U3422 ( .A1(n3562), .A2(n2887), .B1(n2886), .B2(n396), .ZN(n2320)
         );
  OAI22_X1 U3423 ( .A1(n446), .A2(n2891), .B1(n2890), .B2(n396), .ZN(n2324) );
  OAI22_X1 U3424 ( .A1(n446), .A2(n2882), .B1(n2881), .B2(n396), .ZN(n2315) );
  OAI22_X1 U3425 ( .A1(n3461), .A2(n3280), .B1(n2799), .B2(n405), .ZN(n2064)
         );
  OAI22_X1 U3426 ( .A1(n3461), .A2(n2767), .B1(n405), .B2(n3280), .ZN(n2197)
         );
  OAI22_X1 U3427 ( .A1(n434), .A2(n3016), .B1(n3015), .B2(n3642), .ZN(n2453)
         );
  OAI22_X1 U3428 ( .A1(n434), .A2(n2999), .B1(n2998), .B2(n3642), .ZN(n2436)
         );
  OAI22_X1 U3429 ( .A1(n434), .A2(n3023), .B1(n3022), .B2(n3642), .ZN(n2460)
         );
  OAI22_X1 U3430 ( .A1(n434), .A2(n3000), .B1(n2999), .B2(n3642), .ZN(n2437)
         );
  OAI22_X1 U3431 ( .A1(n434), .A2(n3014), .B1(n3013), .B2(n3642), .ZN(n2451)
         );
  OAI22_X1 U3432 ( .A1(n434), .A2(n3024), .B1(n3023), .B2(n3642), .ZN(n2461)
         );
  OAI22_X1 U3433 ( .A1(n434), .A2(n3027), .B1(n3026), .B2(n3642), .ZN(n2464)
         );
  OAI22_X1 U3434 ( .A1(n434), .A2(n3013), .B1(n3012), .B2(n3642), .ZN(n2450)
         );
  OAI22_X1 U3435 ( .A1(n434), .A2(n3002), .B1(n3001), .B2(n3642), .ZN(n2439)
         );
  OAI22_X1 U3436 ( .A1(n434), .A2(n3003), .B1(n3002), .B2(n3642), .ZN(n2440)
         );
  OAI22_X1 U3437 ( .A1(n434), .A2(n3026), .B1(n3025), .B2(n3642), .ZN(n2463)
         );
  OAI22_X1 U3438 ( .A1(n434), .A2(n3022), .B1(n3021), .B2(n3642), .ZN(n2459)
         );
  OAI22_X1 U3439 ( .A1(n434), .A2(n3012), .B1(n3011), .B2(n3642), .ZN(n2449)
         );
  OAI22_X1 U3440 ( .A1(n434), .A2(n3015), .B1(n3014), .B2(n3642), .ZN(n2452)
         );
  OAI22_X1 U3441 ( .A1(n434), .A2(n3006), .B1(n3005), .B2(n3642), .ZN(n2443)
         );
  OAI22_X1 U3442 ( .A1(n3559), .A2(n3056), .B1(n3055), .B2(n381), .ZN(n2494)
         );
  OAI22_X1 U3443 ( .A1(n3559), .A2(n3062), .B1(n3061), .B2(n381), .ZN(n2500)
         );
  OAI22_X1 U3444 ( .A1(n3559), .A2(n3050), .B1(n3049), .B2(n381), .ZN(n2488)
         );
  OAI22_X1 U3445 ( .A1(n3559), .A2(n3054), .B1(n3053), .B2(n381), .ZN(n2492)
         );
  OAI22_X1 U3446 ( .A1(n3559), .A2(n3053), .B1(n3052), .B2(n381), .ZN(n2491)
         );
  OAI22_X1 U3447 ( .A1(n3559), .A2(n3033), .B1(n3032), .B2(n381), .ZN(n2471)
         );
  XNOR2_X2 U3448 ( .A(n3701), .B(n3290), .ZN(n3511) );
  INV_X4 U3449 ( .A(n3511), .ZN(n3700) );
  INV_X4 U3450 ( .A(n327), .ZN(n3290) );
  OAI21_X2 U3451 ( .B1(n785), .B2(n765), .A(n766), .ZN(n3581) );
  INV_X4 U3452 ( .A(n3502), .ZN(n3512) );
  INV_X2 U3453 ( .A(n3512), .ZN(n3513) );
  AND2_X2 U3454 ( .A1(n3241), .A2(n375), .ZN(n3705) );
  XNOR2_X1 U3455 ( .A(n779), .B(n558), .ZN(product[37]) );
  INV_X2 U3456 ( .A(n3623), .ZN(n3625) );
  NOR2_X1 U3457 ( .A1(n1403), .A2(n1430), .ZN(n3514) );
  NOR2_X1 U3458 ( .A1(n1403), .A2(n1430), .ZN(n772) );
  NOR2_X1 U3459 ( .A1(n759), .A2(n754), .ZN(n752) );
  XOR2_X1 U3460 ( .A(n1613), .B(n1586), .Z(n3515) );
  NAND2_X1 U3461 ( .A1(n1584), .A2(n1613), .ZN(n3516) );
  NAND2_X1 U3462 ( .A1(n1584), .A2(n1586), .ZN(n3517) );
  NAND2_X1 U3463 ( .A1(n1613), .A2(n1586), .ZN(n3518) );
  NAND3_X1 U3464 ( .A1(n3516), .A2(n3518), .A3(n3517), .ZN(n1581) );
  NAND2_X2 U3465 ( .A1(n1582), .A2(n1611), .ZN(n804) );
  NAND2_X4 U3466 ( .A1(n3241), .A2(n375), .ZN(n3519) );
  NOR2_X1 U3467 ( .A1(n772), .A2(n3528), .ZN(n3520) );
  NOR2_X1 U3468 ( .A1(n3463), .A2(n3514), .ZN(n767) );
  XNOR2_X1 U3469 ( .A(n3755), .B(n3466), .ZN(n3521) );
  BUF_X1 U3470 ( .A(n773), .Z(n3522) );
  XOR2_X1 U3471 ( .A(n1799), .B(n1778), .Z(n3523) );
  XOR2_X1 U3472 ( .A(n1776), .B(n3523), .Z(n1774) );
  NAND2_X1 U3473 ( .A1(n1776), .A2(n1799), .ZN(n3524) );
  NAND2_X1 U3474 ( .A1(n1776), .A2(n1778), .ZN(n3525) );
  NAND2_X1 U3475 ( .A1(n1799), .A2(n1778), .ZN(n3526) );
  NAND3_X1 U3476 ( .A1(n3524), .A2(n3526), .A3(n3525), .ZN(n1773) );
  AOI21_X1 U3477 ( .B1(n683), .B2(n631), .A(n632), .ZN(n3527) );
  NOR2_X1 U3478 ( .A1(n1774), .A2(n1797), .ZN(n846) );
  AOI21_X1 U3479 ( .B1(n683), .B2(n631), .A(n632), .ZN(n630) );
  NOR2_X1 U3480 ( .A1(n1402), .A2(n3464), .ZN(n3528) );
  INV_X2 U3481 ( .A(n3623), .ZN(n3626) );
  AOI21_X1 U3482 ( .B1(n841), .B2(n837), .A(n838), .ZN(n836) );
  INV_X1 U3483 ( .A(n840), .ZN(n838) );
  NAND2_X1 U3484 ( .A1(n3546), .A2(n770), .ZN(n556) );
  OR2_X4 U3485 ( .A1(n3529), .A2(a[0]), .ZN(n419) );
  XNOR2_X1 U3486 ( .A(n3530), .B(n1553), .ZN(n1551) );
  XNOR2_X1 U3487 ( .A(n1583), .B(n1555), .ZN(n3530) );
  AOI21_X1 U3488 ( .B1(n687), .B2(n673), .A(n676), .ZN(n672) );
  OAI22_X1 U3489 ( .A1(n3562), .A2(n2872), .B1(n2871), .B2(n396), .ZN(n2305)
         );
  OAI22_X1 U3490 ( .A1(n3562), .A2(n2878), .B1(n2877), .B2(n396), .ZN(n2311)
         );
  OAI22_X1 U3491 ( .A1(n3561), .A2(n2866), .B1(n396), .B2(n3283), .ZN(n2299)
         );
  OAI22_X1 U3492 ( .A1(n3562), .A2(n2875), .B1(n2874), .B2(n396), .ZN(n2308)
         );
  OAI22_X1 U3493 ( .A1(n3561), .A2(n2894), .B1(n2893), .B2(n396), .ZN(n2327)
         );
  OAI22_X1 U3494 ( .A1(n3561), .A2(n2869), .B1(n2868), .B2(n396), .ZN(n2302)
         );
  OAI22_X1 U3495 ( .A1(n3561), .A2(n2893), .B1(n2892), .B2(n396), .ZN(n2326)
         );
  OAI22_X1 U3496 ( .A1(n3561), .A2(n2870), .B1(n2869), .B2(n396), .ZN(n2303)
         );
  OAI22_X1 U3497 ( .A1(n3561), .A2(n2895), .B1(n2894), .B2(n396), .ZN(n2328)
         );
  OAI22_X1 U3498 ( .A1(n3561), .A2(n2886), .B1(n2885), .B2(n396), .ZN(n2319)
         );
  OAI22_X1 U3499 ( .A1(n3561), .A2(n2897), .B1(n2896), .B2(n396), .ZN(n2330)
         );
  OAI22_X1 U3500 ( .A1(n446), .A2(n3283), .B1(n2898), .B2(n396), .ZN(n2067) );
  OAI22_X1 U3501 ( .A1(n3562), .A2(n2881), .B1(n2880), .B2(n396), .ZN(n2314)
         );
  OAI22_X1 U3502 ( .A1(n3561), .A2(n2868), .B1(n2867), .B2(n396), .ZN(n2301)
         );
  OAI22_X1 U3503 ( .A1(n3561), .A2(n2871), .B1(n2870), .B2(n396), .ZN(n2304)
         );
  XOR2_X1 U3504 ( .A(n1475), .B(n1502), .Z(n3531) );
  XOR2_X1 U3505 ( .A(n3531), .B(n1500), .Z(n1467) );
  XOR2_X1 U3506 ( .A(n1496), .B(n1469), .Z(n3532) );
  XOR2_X1 U3507 ( .A(n3532), .B(n1467), .Z(n1463) );
  NAND2_X1 U3508 ( .A1(n1475), .A2(n1502), .ZN(n3533) );
  NAND2_X1 U3509 ( .A1(n1475), .A2(n1500), .ZN(n3534) );
  NAND2_X1 U3510 ( .A1(n1502), .A2(n1500), .ZN(n3535) );
  NAND3_X1 U3511 ( .A1(n3533), .A2(n3534), .A3(n3535), .ZN(n1466) );
  NAND2_X1 U3512 ( .A1(n1496), .A2(n1469), .ZN(n3536) );
  NAND2_X1 U3513 ( .A1(n1496), .A2(n1467), .ZN(n3537) );
  NAND2_X1 U3514 ( .A1(n1469), .A2(n1467), .ZN(n3538) );
  NAND3_X1 U3515 ( .A1(n3536), .A2(n3537), .A3(n3538), .ZN(n1462) );
  XOR2_X1 U3516 ( .A(n2506), .B(n2442), .Z(n3539) );
  XOR2_X1 U3517 ( .A(n2538), .B(n3539), .Z(n1509) );
  NAND2_X1 U3518 ( .A1(n2538), .A2(n2506), .ZN(n3540) );
  NAND2_X1 U3519 ( .A1(n2538), .A2(n2442), .ZN(n3541) );
  NAND2_X1 U3520 ( .A1(n2506), .A2(n2442), .ZN(n3542) );
  NAND3_X1 U3521 ( .A1(n3540), .A2(n3542), .A3(n3541), .ZN(n1508) );
  INV_X8 U3522 ( .A(n3543), .ZN(n434) );
  INV_X2 U3523 ( .A(n3426), .ZN(n3640) );
  OAI22_X1 U3524 ( .A1(n434), .A2(n3007), .B1(n3006), .B2(n3641), .ZN(n2444)
         );
  AOI21_X2 U3525 ( .B1(n691), .B2(n615), .A(n616), .ZN(n614) );
  INV_X4 U3526 ( .A(n345), .ZN(n3681) );
  BUF_X1 U3527 ( .A(n3606), .Z(n3545) );
  XOR2_X1 U3528 ( .A(a[28]), .B(n363), .Z(n3229) );
  OR2_X1 U3529 ( .A1(n3464), .A2(n1402), .ZN(n3546) );
  AND2_X2 U3530 ( .A1(n3651), .A2(n3652), .ZN(n808) );
  INV_X4 U3531 ( .A(a[18]), .ZN(n3680) );
  NOR2_X1 U3532 ( .A1(n811), .A2(n814), .ZN(n3547) );
  BUF_X1 U3533 ( .A(n749), .Z(n3548) );
  NAND2_X1 U3534 ( .A1(n1551), .A2(n1581), .ZN(n801) );
  NAND2_X1 U3535 ( .A1(n1011), .A2(n815), .ZN(n565) );
  NAND2_X2 U3536 ( .A1(n3760), .A2(n348), .ZN(n3612) );
  BUF_X1 U3537 ( .A(n1403), .Z(n3549) );
  AOI21_X1 U3538 ( .B1(n761), .B2(n725), .A(n726), .ZN(n3550) );
  AOI21_X1 U3539 ( .B1(n761), .B2(n725), .A(n726), .ZN(n724) );
  NAND2_X4 U3540 ( .A1(n3232), .A2(n3468), .ZN(n3551) );
  NAND2_X4 U3541 ( .A1(n3232), .A2(n3468), .ZN(n3552) );
  OAI22_X1 U3542 ( .A1(n458), .A2(n2759), .B1(n2758), .B2(n3639), .ZN(n2188)
         );
  INV_X1 U3543 ( .A(n324), .ZN(n3291) );
  OAI21_X1 U3544 ( .B1(n800), .B2(n804), .A(n801), .ZN(n3553) );
  INV_X1 U3545 ( .A(n422), .ZN(n3554) );
  INV_X2 U3546 ( .A(n3554), .ZN(n3555) );
  OAI21_X1 U3547 ( .B1(n800), .B2(n804), .A(n801), .ZN(n799) );
  INV_X1 U3548 ( .A(n811), .ZN(n1010) );
  NOR2_X1 U3549 ( .A1(n819), .A2(n824), .ZN(n817) );
  INV_X1 U3550 ( .A(n824), .ZN(n822) );
  OAI22_X1 U3551 ( .A1(n434), .A2(n3005), .B1(n3004), .B2(n3641), .ZN(n2442)
         );
  OAI22_X1 U3552 ( .A1(n3559), .A2(n3044), .B1(n3043), .B2(n381), .ZN(n2482)
         );
  OAI22_X1 U3553 ( .A1(n3559), .A2(n3043), .B1(n3042), .B2(n381), .ZN(n2481)
         );
  OAI22_X1 U3554 ( .A1(n431), .A2(n3046), .B1(n3045), .B2(n381), .ZN(n2484) );
  OAI22_X1 U3555 ( .A1(n431), .A2(n3031), .B1(n381), .B2(n3288), .ZN(n2469) );
  OAI22_X1 U3556 ( .A1(n431), .A2(n3035), .B1(n3034), .B2(n381), .ZN(n2473) );
  OAI22_X1 U3557 ( .A1(n431), .A2(n3039), .B1(n3038), .B2(n381), .ZN(n2477) );
  OAI22_X1 U3558 ( .A1(n431), .A2(n3041), .B1(n3040), .B2(n381), .ZN(n2479) );
  OAI22_X1 U3559 ( .A1(n3579), .A2(n2959), .B1(n2958), .B2(n3650), .ZN(n2394)
         );
  OAI22_X1 U3560 ( .A1(n440), .A2(n2963), .B1(n2962), .B2(n3649), .ZN(n2398)
         );
  OAI22_X1 U3561 ( .A1(n3579), .A2(n2961), .B1(n2960), .B2(n3649), .ZN(n2396)
         );
  OAI22_X1 U3562 ( .A1(n440), .A2(n2936), .B1(n2935), .B2(n3649), .ZN(n2371)
         );
  OAI22_X1 U3563 ( .A1(n3579), .A2(n2935), .B1(n2934), .B2(n3649), .ZN(n2370)
         );
  OAI22_X1 U3564 ( .A1(n440), .A2(n2957), .B1(n2956), .B2(n3649), .ZN(n2392)
         );
  OAI22_X1 U3565 ( .A1(n440), .A2(n2934), .B1(n2933), .B2(n3649), .ZN(n2369)
         );
  OAI22_X1 U3566 ( .A1(n3580), .A2(n2939), .B1(n2938), .B2(n3649), .ZN(n2374)
         );
  OAI22_X1 U3567 ( .A1(n3579), .A2(n2956), .B1(n2955), .B2(n3649), .ZN(n2391)
         );
  OAI22_X1 U3568 ( .A1(n3580), .A2(n2953), .B1(n2952), .B2(n3649), .ZN(n2388)
         );
  OAI22_X1 U3569 ( .A1(n3579), .A2(n2946), .B1(n2945), .B2(n3649), .ZN(n2381)
         );
  OAI22_X1 U3570 ( .A1(n3580), .A2(n2943), .B1(n2942), .B2(n3649), .ZN(n2378)
         );
  OAI22_X1 U3571 ( .A1(n3579), .A2(n2954), .B1(n2953), .B2(n3650), .ZN(n2389)
         );
  OAI22_X1 U3572 ( .A1(n3579), .A2(n2950), .B1(n2949), .B2(n3650), .ZN(n2385)
         );
  OAI22_X1 U3573 ( .A1(n3580), .A2(n2947), .B1(n2946), .B2(n3650), .ZN(n2382)
         );
  OAI22_X1 U3574 ( .A1(n464), .A2(n2673), .B1(n2672), .B2(n3625), .ZN(n2100)
         );
  OAI22_X1 U3575 ( .A1(n464), .A2(n2675), .B1(n2674), .B2(n3626), .ZN(n2102)
         );
  OAI22_X1 U3576 ( .A1(n464), .A2(n2681), .B1(n2680), .B2(n3625), .ZN(n2108)
         );
  OAI22_X1 U3577 ( .A1(n464), .A2(n2676), .B1(n2675), .B2(n3625), .ZN(n2103)
         );
  OAI22_X1 U3578 ( .A1(n464), .A2(n2690), .B1(n2689), .B2(n3626), .ZN(n2117)
         );
  OAI22_X1 U3579 ( .A1(n464), .A2(n2689), .B1(n2688), .B2(n3625), .ZN(n2116)
         );
  OAI22_X1 U3580 ( .A1(n464), .A2(n2680), .B1(n2679), .B2(n3626), .ZN(n2107)
         );
  OAI22_X1 U3581 ( .A1(n464), .A2(n2679), .B1(n2678), .B2(n3626), .ZN(n2106)
         );
  OAI22_X1 U3582 ( .A1(n464), .A2(n2688), .B1(n2687), .B2(n3625), .ZN(n2115)
         );
  OAI22_X1 U3583 ( .A1(n464), .A2(n2692), .B1(n2691), .B2(n3625), .ZN(n2119)
         );
  OAI22_X1 U3584 ( .A1(n464), .A2(n2686), .B1(n2685), .B2(n3625), .ZN(n2113)
         );
  OAI22_X1 U3585 ( .A1(n464), .A2(n2685), .B1(n2684), .B2(n3625), .ZN(n2112)
         );
  OAI22_X1 U3586 ( .A1(n464), .A2(n2684), .B1(n2683), .B2(n3626), .ZN(n2111)
         );
  OAI22_X1 U3587 ( .A1(n464), .A2(n2678), .B1(n2677), .B2(n3626), .ZN(n2105)
         );
  OAI22_X1 U3588 ( .A1(n464), .A2(n2683), .B1(n2682), .B2(n3626), .ZN(n2110)
         );
  OAI22_X1 U3589 ( .A1(n464), .A2(n2695), .B1(n2694), .B2(n3625), .ZN(n2122)
         );
  OAI22_X1 U3590 ( .A1(n464), .A2(n2677), .B1(n2676), .B2(n3625), .ZN(n2104)
         );
  OAI22_X1 U3591 ( .A1(n464), .A2(n2687), .B1(n2686), .B2(n3626), .ZN(n2114)
         );
  OAI22_X1 U3592 ( .A1(n464), .A2(n2694), .B1(n2693), .B2(n3625), .ZN(n2121)
         );
  OAI22_X1 U3593 ( .A1(n464), .A2(n2691), .B1(n2690), .B2(n3626), .ZN(n2118)
         );
  OAI22_X1 U3594 ( .A1(n464), .A2(n2682), .B1(n2681), .B2(n3625), .ZN(n2109)
         );
  OAI22_X1 U3595 ( .A1(n464), .A2(n2693), .B1(n2692), .B2(n3626), .ZN(n2120)
         );
  OAI22_X1 U3596 ( .A1(n464), .A2(n2696), .B1(n2695), .B2(n3626), .ZN(n2123)
         );
  OAI22_X1 U3597 ( .A1(n464), .A2(n2697), .B1(n2696), .B2(n3625), .ZN(n2124)
         );
  OAI22_X1 U3598 ( .A1(n464), .A2(n2699), .B1(n2698), .B2(n3626), .ZN(n2126)
         );
  XNOR2_X1 U3599 ( .A(n679), .B(n544), .ZN(product[51]) );
  OAI22_X1 U3600 ( .A1(n449), .A2(n2841), .B1(n2840), .B2(n399), .ZN(n2273) );
  OAI22_X1 U3601 ( .A1(n449), .A2(n2836), .B1(n2835), .B2(n399), .ZN(n2268) );
  OAI22_X1 U3602 ( .A1(n449), .A2(n2834), .B1(n2833), .B2(n399), .ZN(n2266) );
  OAI22_X1 U3603 ( .A1(n449), .A2(n2851), .B1(n2850), .B2(n399), .ZN(n2283) );
  OAI22_X1 U3604 ( .A1(n449), .A2(n2844), .B1(n2843), .B2(n399), .ZN(n2276) );
  OAI22_X1 U3605 ( .A1(n449), .A2(n2840), .B1(n2839), .B2(n399), .ZN(n2272) );
  OAI22_X1 U3606 ( .A1(n449), .A2(n2857), .B1(n2856), .B2(n399), .ZN(n2289) );
  OAI22_X1 U3607 ( .A1(n449), .A2(n2862), .B1(n2861), .B2(n399), .ZN(n2294) );
  OAI22_X1 U3608 ( .A1(n449), .A2(n2855), .B1(n2854), .B2(n399), .ZN(n2287) );
  OAI22_X1 U3609 ( .A1(n449), .A2(n2850), .B1(n2849), .B2(n399), .ZN(n2282) );
  OAI22_X1 U3610 ( .A1(n449), .A2(n2837), .B1(n2836), .B2(n399), .ZN(n2269) );
  OAI22_X1 U3611 ( .A1(n449), .A2(n2845), .B1(n2844), .B2(n399), .ZN(n2277) );
  OAI22_X1 U3612 ( .A1(n449), .A2(n2854), .B1(n2853), .B2(n399), .ZN(n2286) );
  OAI22_X1 U3613 ( .A1(n449), .A2(n2849), .B1(n2848), .B2(n399), .ZN(n2281) );
  OAI22_X1 U3614 ( .A1(n449), .A2(n2848), .B1(n2847), .B2(n399), .ZN(n2280) );
  OAI22_X1 U3615 ( .A1(n449), .A2(n2860), .B1(n2859), .B2(n399), .ZN(n2292) );
  INV_X1 U3616 ( .A(n3488), .ZN(n3557) );
  NAND2_X4 U3617 ( .A1(n3621), .A2(n3622), .ZN(n3757) );
  NOR2_X4 U3618 ( .A1(n1820), .A2(n1841), .ZN(n861) );
  INV_X1 U3619 ( .A(n3639), .ZN(n3558) );
  OAI22_X1 U3620 ( .A1(n3703), .A2(n3084), .B1(n3083), .B2(n3605), .ZN(n2523)
         );
  OAI22_X1 U3621 ( .A1(n3703), .A2(n3069), .B1(n3068), .B2(n3604), .ZN(n2508)
         );
  OAI22_X1 U3622 ( .A1(n3703), .A2(n3090), .B1(n3089), .B2(n3605), .ZN(n2529)
         );
  OAI22_X1 U3623 ( .A1(n3703), .A2(n3094), .B1(n3093), .B2(n3604), .ZN(n2533)
         );
  OAI22_X1 U3624 ( .A1(n3703), .A2(n3095), .B1(n3094), .B2(n3605), .ZN(n2534)
         );
  OAI22_X1 U3625 ( .A1(n3703), .A2(n3667), .B1(n3096), .B2(n3604), .ZN(n2073)
         );
  OAI22_X1 U3626 ( .A1(n3703), .A2(n3085), .B1(n3084), .B2(n3605), .ZN(n2524)
         );
  OAI22_X1 U3627 ( .A1(n3703), .A2(n3082), .B1(n3081), .B2(n3605), .ZN(n2521)
         );
  OAI22_X1 U3628 ( .A1(n3703), .A2(n3089), .B1(n3088), .B2(n3604), .ZN(n2528)
         );
  OAI22_X1 U3629 ( .A1(n3703), .A2(n3072), .B1(n3071), .B2(n3604), .ZN(n2511)
         );
  OAI22_X1 U3630 ( .A1(n428), .A2(n3087), .B1(n3086), .B2(n3604), .ZN(n2526)
         );
  OAI22_X1 U3631 ( .A1(n428), .A2(n3073), .B1(n3072), .B2(n3605), .ZN(n2512)
         );
  OAI22_X1 U3632 ( .A1(n3703), .A2(n3076), .B1(n3075), .B2(n3604), .ZN(n2515)
         );
  OAI22_X1 U3633 ( .A1(n428), .A2(n3064), .B1(n3605), .B2(n3667), .ZN(n2503)
         );
  OAI22_X1 U3634 ( .A1(n428), .A2(n3066), .B1(n3065), .B2(n3604), .ZN(n2505)
         );
  OAI22_X1 U3635 ( .A1(n3560), .A2(n3060), .B1(n3059), .B2(n381), .ZN(n2498)
         );
  OAI22_X1 U3636 ( .A1(n3560), .A2(n3048), .B1(n3047), .B2(n381), .ZN(n2486)
         );
  OAI22_X1 U3637 ( .A1(n3560), .A2(n3288), .B1(n3063), .B2(n381), .ZN(n2072)
         );
  OAI22_X1 U3638 ( .A1(n3559), .A2(n3061), .B1(n3060), .B2(n381), .ZN(n2499)
         );
  OAI22_X1 U3639 ( .A1(n3559), .A2(n3042), .B1(n3041), .B2(n381), .ZN(n2480)
         );
  OAI22_X1 U3640 ( .A1(n3560), .A2(n3059), .B1(n3058), .B2(n381), .ZN(n2497)
         );
  OAI22_X1 U3641 ( .A1(n3560), .A2(n3052), .B1(n3051), .B2(n381), .ZN(n2490)
         );
  OAI22_X1 U3642 ( .A1(n3560), .A2(n3051), .B1(n3050), .B2(n381), .ZN(n2489)
         );
  OAI22_X1 U3643 ( .A1(n3559), .A2(n3058), .B1(n3057), .B2(n381), .ZN(n2496)
         );
  OAI22_X1 U3644 ( .A1(n3559), .A2(n3045), .B1(n3044), .B2(n381), .ZN(n2483)
         );
  OAI22_X1 U3645 ( .A1(n3560), .A2(n3037), .B1(n3036), .B2(n381), .ZN(n2475)
         );
  OAI22_X1 U3646 ( .A1(n3559), .A2(n3032), .B1(n3031), .B2(n381), .ZN(n2470)
         );
  OAI22_X1 U3647 ( .A1(n3560), .A2(n3049), .B1(n3048), .B2(n381), .ZN(n2487)
         );
  OAI22_X1 U3648 ( .A1(n431), .A2(n3040), .B1(n3039), .B2(n381), .ZN(n2478) );
  OAI22_X1 U3649 ( .A1(n3559), .A2(n3047), .B1(n3046), .B2(n381), .ZN(n2485)
         );
  INV_X2 U3650 ( .A(n3679), .ZN(n3560) );
  INV_X2 U3651 ( .A(n3679), .ZN(n3559) );
  INV_X1 U3652 ( .A(n3679), .ZN(n431) );
  OAI22_X1 U3653 ( .A1(n3456), .A2(n2702), .B1(n2701), .B2(n411), .ZN(n2130)
         );
  OAI22_X1 U3654 ( .A1(n3456), .A2(n2705), .B1(n2704), .B2(n411), .ZN(n2133)
         );
  OAI22_X1 U3655 ( .A1(n3456), .A2(n2704), .B1(n2703), .B2(n411), .ZN(n2132)
         );
  OAI22_X1 U3656 ( .A1(n3456), .A2(n2706), .B1(n2705), .B2(n411), .ZN(n2134)
         );
  OAI22_X1 U3657 ( .A1(n461), .A2(n2712), .B1(n2711), .B2(n411), .ZN(n2140) );
  OAI22_X1 U3658 ( .A1(n3456), .A2(n2707), .B1(n2706), .B2(n411), .ZN(n2135)
         );
  OAI22_X1 U3659 ( .A1(n461), .A2(n2719), .B1(n2718), .B2(n411), .ZN(n2147) );
  OAI22_X1 U3660 ( .A1(n461), .A2(n2717), .B1(n2716), .B2(n411), .ZN(n2145) );
  OAI22_X1 U3661 ( .A1(n461), .A2(n2720), .B1(n2719), .B2(n411), .ZN(n2148) );
  OAI22_X1 U3662 ( .A1(n461), .A2(n2715), .B1(n2714), .B2(n411), .ZN(n2143) );
  OAI22_X1 U3663 ( .A1(n461), .A2(n2723), .B1(n2722), .B2(n411), .ZN(n2151) );
  OAI22_X1 U3664 ( .A1(n461), .A2(n2730), .B1(n2729), .B2(n411), .ZN(n2158) );
  OAI22_X1 U3665 ( .A1(n3456), .A2(n2716), .B1(n2715), .B2(n411), .ZN(n2144)
         );
  OAI22_X1 U3666 ( .A1(n461), .A2(n2727), .B1(n2726), .B2(n411), .ZN(n2155) );
  OAI22_X1 U3667 ( .A1(n461), .A2(n2722), .B1(n2721), .B2(n411), .ZN(n2150) );
  OAI22_X1 U3668 ( .A1(n3660), .A2(n2731), .B1(n2730), .B2(n411), .ZN(n2159)
         );
  XOR2_X2 U3669 ( .A(n1525), .B(n1556), .Z(n3590) );
  XNOR2_X2 U3670 ( .A(n3777), .B(n3490), .ZN(n3689) );
  INV_X2 U3671 ( .A(n3764), .ZN(n3562) );
  INV_X4 U3672 ( .A(n3764), .ZN(n3561) );
  INV_X2 U3673 ( .A(n3563), .ZN(n3564) );
  INV_X1 U3674 ( .A(n3764), .ZN(n446) );
  OR2_X2 U3675 ( .A1(n3712), .A2(n3713), .ZN(n2537) );
  NOR2_X2 U3676 ( .A1(n1489), .A2(n1518), .ZN(n788) );
  NAND2_X2 U3677 ( .A1(n3758), .A2(n336), .ZN(n3621) );
  OAI22_X1 U3678 ( .A1(n446), .A2(n2880), .B1(n2879), .B2(n396), .ZN(n2313) );
  FA_X1 U3679 ( .A(n1493), .B(n1520), .CI(n1491), .S(n3565) );
  OAI21_X1 U3680 ( .B1(n843), .B2(n830), .A(n831), .ZN(n829) );
  INV_X1 U3681 ( .A(n3780), .ZN(n3566) );
  NOR2_X2 U3682 ( .A1(n830), .A2(n842), .ZN(n828) );
  INV_X1 U3683 ( .A(n3291), .ZN(n3778) );
  XOR2_X1 U3684 ( .A(n1529), .B(n1558), .Z(n3567) );
  XOR2_X1 U3685 ( .A(n3567), .B(n1527), .Z(n1523) );
  NAND2_X1 U3686 ( .A1(n1562), .A2(n1537), .ZN(n3568) );
  NAND2_X1 U3687 ( .A1(n1562), .A2(n1535), .ZN(n3569) );
  NAND2_X1 U3688 ( .A1(n1537), .A2(n1535), .ZN(n3570) );
  NAND3_X1 U3689 ( .A1(n3568), .A2(n3569), .A3(n3570), .ZN(n1526) );
  NAND2_X1 U3690 ( .A1(n1529), .A2(n1558), .ZN(n3571) );
  NAND2_X1 U3691 ( .A1(n1529), .A2(n1527), .ZN(n3572) );
  NAND2_X1 U3692 ( .A1(n1558), .A2(n1527), .ZN(n3573) );
  NAND3_X1 U3693 ( .A1(n3571), .A2(n3572), .A3(n3573), .ZN(n1522) );
  NOR2_X2 U3694 ( .A1(n1458), .A2(n1431), .ZN(n777) );
  OAI21_X1 U3695 ( .B1(n682), .B2(n680), .A(n681), .ZN(n679) );
  INV_X1 U3696 ( .A(n3738), .ZN(n414) );
  XOR2_X1 U3697 ( .A(n1751), .B(n1728), .Z(n3574) );
  XOR2_X1 U3698 ( .A(n1726), .B(n3574), .Z(n1724) );
  NAND2_X1 U3699 ( .A1(n1726), .A2(n1751), .ZN(n3575) );
  NAND2_X1 U3700 ( .A1(n1726), .A2(n1728), .ZN(n3576) );
  NAND2_X1 U3701 ( .A1(n1751), .A2(n1728), .ZN(n3577) );
  NAND3_X1 U3702 ( .A1(n3575), .A2(n3577), .A3(n3576), .ZN(n1723) );
  BUF_X1 U3703 ( .A(n761), .Z(n3578) );
  NOR2_X1 U3704 ( .A1(n1698), .A2(n1723), .ZN(n824) );
  AND2_X4 U3705 ( .A1(n3236), .A2(n3648), .ZN(n3688) );
  OAI21_X1 U3706 ( .B1(n785), .B2(n765), .A(n766), .ZN(n764) );
  OAI22_X1 U3707 ( .A1(n464), .A2(n3500), .B1(n2700), .B2(n3625), .ZN(n2061)
         );
  OAI21_X2 U3708 ( .B1(n531), .B2(n604), .A(n605), .ZN(n603) );
  OAI22_X1 U3709 ( .A1(n3561), .A2(n2884), .B1(n2883), .B2(n396), .ZN(n2317)
         );
  OAI21_X1 U3710 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  OAI22_X1 U3711 ( .A1(n3579), .A2(n2952), .B1(n2951), .B2(n3650), .ZN(n2387)
         );
  INV_X2 U3712 ( .A(n3705), .ZN(n425) );
  OAI21_X1 U3713 ( .B1(n744), .B2(n3458), .A(n739), .ZN(n737) );
  OAI22_X1 U3714 ( .A1(n3562), .A2(n2896), .B1(n2895), .B2(n396), .ZN(n2329)
         );
  BUF_X1 U3715 ( .A(n706), .Z(n3582) );
  INV_X2 U3716 ( .A(n321), .ZN(n3583) );
  INV_X1 U3717 ( .A(n321), .ZN(n3292) );
  OAI22_X1 U3718 ( .A1(n458), .A2(n2761), .B1(n2760), .B2(n3638), .ZN(n2190)
         );
  INV_X4 U3719 ( .A(a[30]), .ZN(n3739) );
  NAND2_X1 U3720 ( .A1(n3584), .A2(n3585), .ZN(n3587) );
  INV_X1 U3721 ( .A(n3629), .ZN(n3584) );
  INV_X2 U3722 ( .A(n3585), .ZN(n3588) );
  OR2_X4 U3723 ( .A1(n3589), .A2(n3704), .ZN(n455) );
  INV_X8 U3724 ( .A(n3704), .ZN(n405) );
  NAND2_X2 U3725 ( .A1(n1351), .A2(n1376), .ZN(n760) );
  NOR2_X2 U3726 ( .A1(n1670), .A2(n1697), .ZN(n819) );
  NAND2_X1 U3727 ( .A1(n1670), .A2(n1697), .ZN(n820) );
  OAI22_X1 U3728 ( .A1(n419), .A2(n3292), .B1(n3195), .B2(n369), .ZN(n2076) );
  OAI22_X1 U3729 ( .A1(n419), .A2(n3163), .B1(n3292), .B2(n369), .ZN(n2605) );
  NAND2_X1 U3730 ( .A1(n995), .A2(n716), .ZN(n549) );
  INV_X1 U3731 ( .A(n686), .ZN(n684) );
  NAND2_X1 U3732 ( .A1(n686), .A2(n673), .ZN(n671) );
  AOI21_X2 U3733 ( .B1(n995), .B2(n721), .A(n714), .ZN(n712) );
  NAND2_X2 U3734 ( .A1(n996), .A2(n995), .ZN(n711) );
  INV_X1 U3735 ( .A(n3705), .ZN(n3698) );
  OAI22_X1 U3736 ( .A1(n3703), .A2(n3091), .B1(n3090), .B2(n3604), .ZN(n2530)
         );
  OAI22_X1 U3737 ( .A1(n3703), .A2(n3079), .B1(n3078), .B2(n3605), .ZN(n2518)
         );
  OAI22_X1 U3738 ( .A1(n3703), .A2(n3093), .B1(n3092), .B2(n3604), .ZN(n2532)
         );
  OAI22_X1 U3739 ( .A1(n3703), .A2(n3075), .B1(n3074), .B2(n3605), .ZN(n2514)
         );
  OAI22_X1 U3740 ( .A1(n3703), .A2(n3092), .B1(n3091), .B2(n3605), .ZN(n2531)
         );
  OAI22_X1 U3741 ( .A1(n3703), .A2(n3088), .B1(n3087), .B2(n3604), .ZN(n2527)
         );
  OAI22_X1 U3742 ( .A1(n3703), .A2(n3086), .B1(n3085), .B2(n3604), .ZN(n2525)
         );
  OAI22_X1 U3743 ( .A1(n3703), .A2(n3083), .B1(n3082), .B2(n3604), .ZN(n2522)
         );
  OAI22_X1 U3744 ( .A1(n3703), .A2(n3078), .B1(n3077), .B2(n3605), .ZN(n2517)
         );
  OAI22_X1 U3745 ( .A1(n3703), .A2(n3074), .B1(n3073), .B2(n3605), .ZN(n2513)
         );
  OAI22_X1 U3746 ( .A1(n428), .A2(n3081), .B1(n3080), .B2(n3605), .ZN(n2520)
         );
  OAI22_X1 U3747 ( .A1(n3703), .A2(n3070), .B1(n3069), .B2(n3605), .ZN(n2509)
         );
  OAI22_X1 U3748 ( .A1(n428), .A2(n3077), .B1(n3076), .B2(n3605), .ZN(n2516)
         );
  OAI22_X1 U3749 ( .A1(n428), .A2(n3080), .B1(n3079), .B2(n3604), .ZN(n2519)
         );
  OAI22_X1 U3750 ( .A1(n428), .A2(n3065), .B1(n3064), .B2(n3605), .ZN(n2504)
         );
  XOR2_X2 U3751 ( .A(n3590), .B(n1554), .Z(n1521) );
  NAND2_X1 U3752 ( .A1(n1525), .A2(n1556), .ZN(n3591) );
  NAND2_X1 U3753 ( .A1(n1525), .A2(n1554), .ZN(n3592) );
  NAND2_X1 U3754 ( .A1(n1556), .A2(n1554), .ZN(n3593) );
  NAND3_X1 U3755 ( .A1(n3591), .A2(n3592), .A3(n3593), .ZN(n1520) );
  NAND2_X1 U3756 ( .A1(n1552), .A2(n1523), .ZN(n3594) );
  NAND2_X1 U3757 ( .A1(n1552), .A2(n1521), .ZN(n3595) );
  NAND2_X1 U3758 ( .A1(n1523), .A2(n1521), .ZN(n3596) );
  NAND3_X2 U3759 ( .A1(n3594), .A2(n3595), .A3(n3596), .ZN(n1518) );
  NAND2_X1 U3760 ( .A1(n753), .A2(n729), .ZN(n3597) );
  INV_X1 U3761 ( .A(n730), .ZN(n3598) );
  AND2_X2 U3762 ( .A1(n3597), .A2(n3598), .ZN(n728) );
  INV_X1 U3763 ( .A(n3469), .ZN(n3599) );
  NOR2_X2 U3764 ( .A1(n731), .A2(n747), .ZN(n729) );
  XNOR2_X1 U3765 ( .A(n2542), .B(n3600), .ZN(n1636) );
  XNOR2_X2 U3766 ( .A(n2318), .B(n2510), .ZN(n3600) );
  XNOR2_X1 U3767 ( .A(n717), .B(n549), .ZN(product[46]) );
  INV_X16 U3768 ( .A(n465), .ZN(n3784) );
  XNOR2_X1 U3769 ( .A(n3737), .B(n3583), .ZN(n3601) );
  OAI21_X1 U3770 ( .B1(n724), .B2(n718), .A(n719), .ZN(n717) );
  OAI22_X1 U3771 ( .A1(n422), .A2(n3143), .B1(n3142), .B2(n372), .ZN(n2584) );
  NAND2_X1 U3772 ( .A1(n1820), .A2(n1841), .ZN(n862) );
  INV_X4 U3773 ( .A(n3511), .ZN(n3602) );
  INV_X1 U3774 ( .A(n3602), .ZN(n3603) );
  INV_X4 U3775 ( .A(n3602), .ZN(n3605) );
  INV_X4 U3776 ( .A(n3602), .ZN(n3604) );
  INV_X1 U3777 ( .A(n794), .ZN(n792) );
  NOR2_X2 U3778 ( .A1(n3565), .A2(n1518), .ZN(n3606) );
  NAND2_X1 U3779 ( .A1(n3781), .A2(n342), .ZN(n3609) );
  NAND2_X1 U3780 ( .A1(n3607), .A2(n3608), .ZN(n3610) );
  NAND2_X1 U3781 ( .A1(n3609), .A2(n3610), .ZN(n3780) );
  INV_X1 U3782 ( .A(n3781), .ZN(n3607) );
  INV_X1 U3783 ( .A(n3780), .ZN(n393) );
  NAND2_X1 U3784 ( .A1(n3611), .A2(n3644), .ZN(n3613) );
  NAND2_X2 U3785 ( .A1(n3612), .A2(n3613), .ZN(n3759) );
  INV_X1 U3786 ( .A(n3760), .ZN(n3611) );
  OAI22_X1 U3787 ( .A1(n449), .A2(n2853), .B1(n2852), .B2(n399), .ZN(n2285) );
  NAND2_X1 U3788 ( .A1(n3614), .A2(n3615), .ZN(n3617) );
  NAND2_X2 U3789 ( .A1(n3616), .A2(n3617), .ZN(n3753) );
  INV_X1 U3790 ( .A(n3754), .ZN(n3614) );
  INV_X1 U3791 ( .A(n360), .ZN(n3615) );
  OAI21_X1 U3792 ( .B1(n3763), .B2(n3700), .A(n330), .ZN(n2502) );
  AOI21_X1 U3793 ( .B1(n806), .B2(n763), .A(n764), .ZN(n3618) );
  NAND2_X1 U3794 ( .A1(n3619), .A2(n3620), .ZN(n3622) );
  INV_X1 U3795 ( .A(n3457), .ZN(n3619) );
  INV_X1 U3796 ( .A(n336), .ZN(n3620) );
  AOI21_X1 U3797 ( .B1(n3485), .B2(n806), .A(n3581), .ZN(n3684) );
  INV_X4 U3798 ( .A(n3657), .ZN(n449) );
  INV_X4 U3799 ( .A(n3657), .ZN(n3643) );
  OAI21_X1 U3800 ( .B1(n3657), .B2(n3759), .A(n3588), .ZN(n2264) );
  OAI21_X1 U3801 ( .B1(n3670), .B2(n3780), .A(n3564), .ZN(n2332) );
  OAI22_X1 U3802 ( .A1(n3456), .A2(n2701), .B1(n411), .B2(n3278), .ZN(n2129)
         );
  OAI22_X1 U3803 ( .A1(n461), .A2(n2703), .B1(n2702), .B2(n411), .ZN(n2131) );
  OAI22_X1 U3804 ( .A1(n461), .A2(n2709), .B1(n2708), .B2(n411), .ZN(n2137) );
  OAI22_X1 U3805 ( .A1(n461), .A2(n2708), .B1(n2707), .B2(n411), .ZN(n2136) );
  OAI22_X1 U3806 ( .A1(n461), .A2(n2721), .B1(n2720), .B2(n411), .ZN(n2149) );
  OAI22_X1 U3807 ( .A1(n3456), .A2(n2711), .B1(n2710), .B2(n411), .ZN(n2139)
         );
  OAI22_X1 U3808 ( .A1(n3456), .A2(n2713), .B1(n2712), .B2(n411), .ZN(n2141)
         );
  OAI22_X1 U3809 ( .A1(n461), .A2(n2710), .B1(n2709), .B2(n411), .ZN(n2138) );
  OAI22_X1 U3810 ( .A1(n461), .A2(n2718), .B1(n2717), .B2(n411), .ZN(n2146) );
  OAI22_X1 U3811 ( .A1(n461), .A2(n2724), .B1(n2723), .B2(n411), .ZN(n2152) );
  OAI22_X1 U3812 ( .A1(n461), .A2(n2725), .B1(n2724), .B2(n411), .ZN(n2153) );
  OAI22_X1 U3813 ( .A1(n461), .A2(n2714), .B1(n2713), .B2(n411), .ZN(n2142) );
  OAI22_X1 U3814 ( .A1(n3456), .A2(n2732), .B1(n2731), .B2(n411), .ZN(n2160)
         );
  OAI22_X1 U3815 ( .A1(n461), .A2(n3278), .B1(n2733), .B2(n411), .ZN(n2062) );
  OAI22_X1 U3816 ( .A1(n461), .A2(n2726), .B1(n2725), .B2(n411), .ZN(n2154) );
  OAI22_X1 U3817 ( .A1(n3660), .A2(n2729), .B1(n2728), .B2(n411), .ZN(n2157)
         );
  OAI22_X1 U3818 ( .A1(n3660), .A2(n2728), .B1(n2727), .B2(n411), .ZN(n2156)
         );
  INV_X2 U3819 ( .A(n414), .ZN(n3623) );
  INV_X1 U3820 ( .A(n3623), .ZN(n3624) );
  XNOR2_X1 U3821 ( .A(n2547), .B(n3627), .ZN(n1768) );
  XNOR2_X1 U3822 ( .A(n2323), .B(n2355), .ZN(n3627) );
  OAI22_X1 U3823 ( .A1(n3416), .A2(n2978), .B1(n2977), .B2(n387), .ZN(n2414)
         );
  INV_X2 U3824 ( .A(n3601), .ZN(n3628) );
  OAI22_X1 U3825 ( .A1(n3551), .A2(n2819), .B1(n2818), .B2(n3469), .ZN(n2250)
         );
  OAI22_X1 U3826 ( .A1(n3551), .A2(n2817), .B1(n2816), .B2(n3468), .ZN(n2248)
         );
  NAND2_X1 U3827 ( .A1(n752), .A2(n729), .ZN(n3630) );
  OR2_X2 U3828 ( .A1(n443), .A2(n2921), .ZN(n3631) );
  OR2_X1 U3829 ( .A1(n2920), .A2(n3656), .ZN(n3632) );
  NAND2_X2 U3830 ( .A1(n3631), .A2(n3632), .ZN(n2355) );
  INV_X2 U3831 ( .A(n3633), .ZN(n3634) );
  XNOR2_X1 U3832 ( .A(n487), .B(n3556), .ZN(n2920) );
  OAI22_X1 U3833 ( .A1(n464), .A2(n2698), .B1(n2697), .B2(n3626), .ZN(n2125)
         );
  INV_X1 U3834 ( .A(n3636), .ZN(n3637) );
  INV_X2 U3835 ( .A(n3640), .ZN(n3642) );
  INV_X4 U3836 ( .A(n3640), .ZN(n3641) );
  OAI21_X1 U3837 ( .B1(n3671), .B2(n3753), .A(n363), .ZN(n2128) );
  INV_X2 U3838 ( .A(n3644), .ZN(n3645) );
  NOR2_X1 U3839 ( .A1(n861), .A2(n864), .ZN(n3646) );
  OAI22_X1 U3840 ( .A1(n3552), .A2(n2823), .B1(n2822), .B2(n3469), .ZN(n2254)
         );
  OAI22_X1 U3841 ( .A1(n3551), .A2(n2821), .B1(n2820), .B2(n3469), .ZN(n2252)
         );
  INV_X2 U3842 ( .A(n390), .ZN(n3647) );
  INV_X1 U3843 ( .A(n752), .ZN(n750) );
  NAND2_X1 U3844 ( .A1(n818), .A2(n809), .ZN(n3651) );
  INV_X1 U3845 ( .A(n810), .ZN(n3652) );
  NAND2_X1 U3846 ( .A1(n1642), .A2(n1669), .ZN(n815) );
  BUF_X1 U3847 ( .A(n464), .Z(n3653) );
  INV_X1 U3848 ( .A(n747), .ZN(n999) );
  NOR2_X2 U3849 ( .A1(n1303), .A2(n1326), .ZN(n747) );
  NAND2_X2 U3850 ( .A1(n1303), .A2(n1326), .ZN(n748) );
  INV_X1 U3851 ( .A(n734), .ZN(n3654) );
  INV_X1 U3852 ( .A(n736), .ZN(n734) );
  NAND2_X1 U3853 ( .A1(n1259), .A2(n1280), .ZN(n736) );
  INV_X1 U3854 ( .A(n738), .ZN(n998) );
  INV_X1 U3855 ( .A(n3659), .ZN(n739) );
  AOI21_X4 U3856 ( .B1(n844), .B2(n852), .A(n845), .ZN(n843) );
  INV_X1 U3857 ( .A(n847), .ZN(n845) );
  INV_X1 U3858 ( .A(n850), .ZN(n852) );
  OAI22_X1 U3859 ( .A1(n3551), .A2(n2830), .B1(n2829), .B2(n3469), .ZN(n2261)
         );
  NOR2_X2 U3860 ( .A1(n1327), .A2(n1350), .ZN(n754) );
  INV_X2 U3861 ( .A(n393), .ZN(n3655) );
  INV_X8 U3862 ( .A(n3655), .ZN(n3656) );
  OAI22_X1 U3863 ( .A1(n458), .A2(n2763), .B1(n2762), .B2(n3639), .ZN(n2192)
         );
  AND2_X1 U3864 ( .A1(n1281), .A2(n1302), .ZN(n3659) );
  OAI22_X1 U3865 ( .A1(n443), .A2(n2914), .B1(n2913), .B2(n3656), .ZN(n2348)
         );
  AND2_X2 U3866 ( .A1(n3233), .A2(n3510), .ZN(n3657) );
  OAI22_X1 U3867 ( .A1(n3551), .A2(n2822), .B1(n2821), .B2(n3469), .ZN(n2253)
         );
  OAI21_X1 U3868 ( .B1(n3635), .B2(n3757), .A(n339), .ZN(n2400) );
  OAI22_X1 U3869 ( .A1(n3643), .A2(n2846), .B1(n2845), .B2(n399), .ZN(n2278)
         );
  OAI22_X1 U3870 ( .A1(n434), .A2(n3019), .B1(n3018), .B2(n3641), .ZN(n2456)
         );
  OAI21_X1 U3871 ( .B1(n3543), .B2(n3751), .A(n336), .ZN(n2434) );
  AOI21_X2 U3872 ( .B1(n3646), .B2(n868), .A(n860), .ZN(n858) );
  BUF_X1 U3873 ( .A(n793), .Z(n3658) );
  OAI22_X1 U3874 ( .A1(n422), .A2(n3132), .B1(n3131), .B2(n372), .ZN(n2573) );
  AND2_X2 U3875 ( .A1(n3230), .A2(n3637), .ZN(n3662) );
  INV_X8 U3876 ( .A(n3662), .ZN(n458) );
  INV_X1 U3877 ( .A(n797), .ZN(n3663) );
  XNOR2_X1 U3878 ( .A(n3664), .B(n1541), .ZN(n1531) );
  XNOR2_X1 U3879 ( .A(n1545), .B(n1543), .ZN(n3664) );
  OAI22_X1 U3880 ( .A1(n3552), .A2(n2818), .B1(n2817), .B2(n3468), .ZN(n2249)
         );
  BUF_X1 U3881 ( .A(n3491), .Z(n3665) );
  NAND2_X2 U3882 ( .A1(n3767), .A2(n330), .ZN(n3668) );
  NAND2_X1 U3883 ( .A1(n3666), .A2(n3667), .ZN(n3669) );
  NAND2_X2 U3884 ( .A1(n3668), .A2(n3669), .ZN(n3766) );
  INV_X1 U3885 ( .A(n3767), .ZN(n3666) );
  AND2_X2 U3886 ( .A1(n3235), .A2(n3566), .ZN(n3670) );
  INV_X8 U3887 ( .A(n3670), .ZN(n443) );
  OAI21_X1 U3888 ( .B1(n3672), .B2(n3628), .A(n3778), .ZN(n2570) );
  NOR2_X2 U3889 ( .A1(n1612), .A2(n1641), .ZN(n811) );
  INV_X1 U3890 ( .A(n835), .ZN(n833) );
  OAI21_X1 U3891 ( .B1(n3661), .B2(n3599), .A(n354), .ZN(n2230) );
  NAND2_X1 U3892 ( .A1(n1123), .A2(n1136), .ZN(n669) );
  NOR2_X1 U3893 ( .A1(n1123), .A2(n1136), .ZN(n668) );
  AOI21_X2 U3894 ( .B1(n658), .B2(n667), .A(n659), .ZN(n657) );
  OAI21_X1 U3895 ( .B1(n657), .B2(n637), .A(n638), .ZN(n636) );
  INV_X1 U3896 ( .A(n657), .ZN(n655) );
  OAI21_X2 U3897 ( .B1(n531), .B2(n684), .A(n685), .ZN(n683) );
  OAI21_X2 U3898 ( .B1(n805), .B2(n784), .A(n3779), .ZN(n783) );
  NAND2_X1 U3899 ( .A1(n1327), .A2(n1350), .ZN(n755) );
  OAI22_X1 U3900 ( .A1(n3552), .A2(n2815), .B1(n2814), .B2(n3468), .ZN(n2246)
         );
  INV_X8 U3901 ( .A(n3672), .ZN(n422) );
  INV_X1 U3902 ( .A(n3658), .ZN(n791) );
  OAI21_X1 U3903 ( .B1(n3662), .B2(n3558), .A(n360), .ZN(n2162) );
  NAND2_X1 U3904 ( .A1(n998), .A2(n739), .ZN(n552) );
  NAND2_X1 U3905 ( .A1(n786), .A2(n799), .ZN(n3673) );
  INV_X1 U3906 ( .A(n787), .ZN(n3674) );
  AND2_X2 U3907 ( .A1(n3673), .A2(n3674), .ZN(n785) );
  NAND2_X1 U3908 ( .A1(a[24]), .A2(n3676), .ZN(n3677) );
  NAND2_X2 U3909 ( .A1(n3675), .A2(n354), .ZN(n3678) );
  INV_X2 U3910 ( .A(a[24]), .ZN(n3675) );
  INV_X2 U3911 ( .A(n354), .ZN(n3676) );
  INV_X8 U3912 ( .A(n3699), .ZN(n396) );
  OAI21_X1 U3913 ( .B1(n3688), .B2(n3471), .A(n3634), .ZN(n2366) );
  NOR2_X1 U3914 ( .A1(n1351), .A2(n1376), .ZN(n759) );
  OAI21_X1 U3915 ( .B1(n3679), .B2(n3766), .A(n333), .ZN(n2468) );
  OAI21_X2 U3916 ( .B1(n754), .B2(n760), .A(n755), .ZN(n753) );
  INV_X1 U3917 ( .A(n3497), .ZN(n1000) );
  NOR2_X1 U3918 ( .A1(n3561), .A2(n2885), .ZN(n3685) );
  NOR2_X1 U3919 ( .A1(n2884), .A2(n396), .ZN(n3686) );
  OR2_X2 U3920 ( .A1(n3685), .A2(n3686), .ZN(n2318) );
  AOI21_X2 U3921 ( .B1(n806), .B2(n3486), .A(n3581), .ZN(n531) );
  XNOR2_X1 U3922 ( .A(n491), .B(n348), .ZN(n2885) );
  OAI21_X1 U3923 ( .B1(n3786), .B2(n3704), .A(n3467), .ZN(n2196) );
  AND2_X2 U3924 ( .A1(n3228), .A2(n3624), .ZN(n3687) );
  INV_X8 U3925 ( .A(n3687), .ZN(n464) );
  OAI22_X1 U3926 ( .A1(n3580), .A2(n2949), .B1(n2948), .B2(n3649), .ZN(n2384)
         );
  OAI21_X1 U3927 ( .B1(n3764), .B2(n3699), .A(n3645), .ZN(n2298) );
  OAI21_X1 U3928 ( .B1(n3687), .B2(n3738), .A(n366), .ZN(n3787) );
  OAI21_X1 U3929 ( .B1(n728), .B2(n613), .A(n614), .ZN(n612) );
  INV_X4 U3930 ( .A(n3689), .ZN(n375) );
  NAND2_X1 U3931 ( .A1(n1009), .A2(n804), .ZN(n563) );
  NOR2_X1 U3932 ( .A1(n1582), .A2(n1611), .ZN(n803) );
  NAND2_X1 U3933 ( .A1(n2542), .A2(n2318), .ZN(n3691) );
  NAND2_X1 U3934 ( .A1(n2542), .A2(n2510), .ZN(n3692) );
  NAND2_X1 U3935 ( .A1(n2318), .A2(n2510), .ZN(n3693) );
  NAND3_X1 U3936 ( .A1(n3691), .A2(n3693), .A3(n3692), .ZN(n1635) );
  BUF_X1 U3937 ( .A(n603), .Z(n3694) );
  OAI22_X1 U3938 ( .A1(n3703), .A2(n3071), .B1(n3070), .B2(n3605), .ZN(n2510)
         );
  INV_X1 U3939 ( .A(n800), .ZN(n1008) );
  OAI21_X1 U3940 ( .B1(n3557), .B2(n3705), .A(n327), .ZN(n2536) );
  NOR2_X2 U3941 ( .A1(n1642), .A2(n1669), .ZN(n814) );
  NAND2_X1 U3942 ( .A1(n1553), .A2(n1583), .ZN(n3695) );
  NAND2_X1 U3943 ( .A1(n1553), .A2(n1555), .ZN(n3696) );
  NAND2_X1 U3944 ( .A1(n1583), .A2(n1555), .ZN(n3697) );
  NAND3_X1 U3945 ( .A1(n3695), .A2(n3697), .A3(n3696), .ZN(n1550) );
  NOR2_X2 U3946 ( .A1(n1551), .A2(n1581), .ZN(n800) );
  NAND2_X1 U3947 ( .A1(n1862), .A2(n1881), .ZN(n870) );
  AOI21_X1 U3948 ( .B1(n826), .B2(n817), .A(n3418), .ZN(n816) );
  NAND2_X2 U3949 ( .A1(n1698), .A2(n1723), .ZN(n825) );
  NAND2_X1 U3950 ( .A1(n1774), .A2(n1797), .ZN(n847) );
  INV_X1 U3951 ( .A(n3504), .ZN(n876) );
  NOR2_X2 U3952 ( .A1(n784), .A2(n765), .ZN(n763) );
  INV_X16 U3953 ( .A(a[0]), .ZN(n369) );
  NAND2_X1 U3954 ( .A1(n844), .A2(n847), .ZN(n570) );
  NAND2_X1 U3955 ( .A1(n844), .A2(n851), .ZN(n842) );
  OAI22_X1 U3956 ( .A1(n3519), .A2(n3116), .B1(n3115), .B2(n3488), .ZN(n2556)
         );
  OAI22_X1 U3957 ( .A1(n3519), .A2(n3128), .B1(n3127), .B2(n3488), .ZN(n2568)
         );
  OAI22_X1 U3958 ( .A1(n3498), .A2(n3125), .B1(n3124), .B2(n3488), .ZN(n2565)
         );
  OAI22_X1 U3959 ( .A1(n425), .A2(n3126), .B1(n3125), .B2(n3488), .ZN(n2566)
         );
  OAI22_X1 U3960 ( .A1(n3519), .A2(n3124), .B1(n3123), .B2(n3488), .ZN(n2564)
         );
  OAI22_X1 U3961 ( .A1(n425), .A2(n3119), .B1(n3118), .B2(n3488), .ZN(n2559)
         );
  OAI22_X1 U3962 ( .A1(n425), .A2(n3122), .B1(n3121), .B2(n3488), .ZN(n2562)
         );
  OAI22_X1 U3963 ( .A1(n3519), .A2(n3117), .B1(n3116), .B2(n3488), .ZN(n2557)
         );
  OAI22_X1 U3964 ( .A1(n3519), .A2(n3120), .B1(n3119), .B2(n3488), .ZN(n2560)
         );
  OAI22_X1 U3965 ( .A1(n3519), .A2(n3118), .B1(n3117), .B2(n3488), .ZN(n2558)
         );
  OAI22_X1 U3966 ( .A1(n3519), .A2(n3111), .B1(n3110), .B2(n375), .ZN(n2551)
         );
  OAI22_X1 U3967 ( .A1(n425), .A2(n3115), .B1(n3114), .B2(n375), .ZN(n2555) );
  OAI22_X1 U3968 ( .A1(n3519), .A2(n3109), .B1(n3108), .B2(n375), .ZN(n2549)
         );
  OAI21_X1 U3969 ( .B1(n866), .B2(n864), .A(n865), .ZN(n863) );
  INV_X1 U3970 ( .A(n864), .ZN(n1019) );
  NAND2_X1 U3971 ( .A1(n859), .A2(n867), .ZN(n857) );
  NOR2_X1 U3972 ( .A1(n861), .A2(n864), .ZN(n859) );
  OAI21_X1 U3973 ( .B1(n816), .B2(n814), .A(n3427), .ZN(n813) );
  INV_X1 U3974 ( .A(n814), .ZN(n1011) );
  NOR2_X1 U3975 ( .A1(n814), .A2(n811), .ZN(n809) );
  OAI22_X1 U3976 ( .A1(n425), .A2(n3103), .B1(n3102), .B2(n375), .ZN(n2543) );
  OAI22_X1 U3977 ( .A1(n3519), .A2(n3098), .B1(n3097), .B2(n3488), .ZN(n2538)
         );
  OAI22_X1 U3978 ( .A1(n425), .A2(n3104), .B1(n3103), .B2(n375), .ZN(n2544) );
  OAI22_X1 U3979 ( .A1(n3519), .A2(n3113), .B1(n3112), .B2(n375), .ZN(n2553)
         );
  OAI22_X1 U3980 ( .A1(n3519), .A2(n3112), .B1(n3111), .B2(n375), .ZN(n2552)
         );
  OAI22_X1 U3981 ( .A1(n3519), .A2(n3099), .B1(n3098), .B2(n375), .ZN(n2539)
         );
  OAI22_X1 U3982 ( .A1(n3519), .A2(n3110), .B1(n3109), .B2(n3488), .ZN(n2550)
         );
  OAI22_X1 U3983 ( .A1(n3519), .A2(n3101), .B1(n3100), .B2(n375), .ZN(n2541)
         );
  NAND2_X1 U3984 ( .A1(n1612), .A2(n1641), .ZN(n812) );
  OAI22_X1 U3985 ( .A1(n3507), .A2(n3121), .B1(n3120), .B2(n3488), .ZN(n2561)
         );
  OAI22_X1 U3986 ( .A1(n3507), .A2(n3438), .B1(n3129), .B2(n3488), .ZN(n2074)
         );
  OAI22_X1 U3987 ( .A1(n3519), .A2(n3127), .B1(n3126), .B2(n3488), .ZN(n2567)
         );
  OAI22_X1 U3988 ( .A1(n3519), .A2(n3123), .B1(n3122), .B2(n3488), .ZN(n2563)
         );
  OAI22_X1 U3989 ( .A1(n3519), .A2(n3105), .B1(n3104), .B2(n3488), .ZN(n2545)
         );
  OAI22_X1 U3990 ( .A1(n425), .A2(n3108), .B1(n3107), .B2(n375), .ZN(n2548) );
  OAI22_X1 U3991 ( .A1(n425), .A2(n3114), .B1(n3113), .B2(n375), .ZN(n2554) );
  OAI22_X1 U3992 ( .A1(n3519), .A2(n3102), .B1(n3101), .B2(n3488), .ZN(n2542)
         );
  OAI22_X1 U3993 ( .A1(n425), .A2(n3106), .B1(n3105), .B2(n375), .ZN(n2546) );
  AOI21_X2 U3994 ( .B1(n670), .B2(n989), .A(n667), .ZN(n665) );
  OAI21_X1 U3995 ( .B1(n3684), .B2(n750), .A(n751), .ZN(n749) );
  OAI21_X1 U3996 ( .B1(n3684), .B2(n707), .A(n708), .ZN(n706) );
  INV_X1 U3997 ( .A(n531), .ZN(n761) );
  NOR2_X2 U3998 ( .A1(n1519), .A2(n1550), .ZN(n793) );
  BUF_X2 U3999 ( .A(n2507), .Z(n3702) );
  INV_X4 U4000 ( .A(n3763), .ZN(n3703) );
  AOI21_X2 U4001 ( .B1(n706), .B2(n994), .A(n703), .ZN(n701) );
  OAI21_X1 U4002 ( .B1(n630), .B2(n624), .A(n625), .ZN(n623) );
  INV_X1 U4003 ( .A(n683), .ZN(n682) );
  NAND2_X1 U4004 ( .A1(n1006), .A2(n789), .ZN(n560) );
  XOR2_X1 U4005 ( .A(n790), .B(n560), .Z(product[35]) );
  NAND2_X1 U4006 ( .A1(n1433), .A2(n1460), .ZN(n3706) );
  NAND2_X1 U4007 ( .A1(n1433), .A2(n1435), .ZN(n3707) );
  NAND2_X1 U4008 ( .A1(n1460), .A2(n1435), .ZN(n3708) );
  NAND3_X1 U4009 ( .A1(n3706), .A2(n3708), .A3(n3707), .ZN(n1430) );
  NOR2_X1 U4010 ( .A1(n1431), .A2(n1458), .ZN(n3709) );
  AOI21_X2 U4011 ( .B1(n856), .B2(n828), .A(n829), .ZN(n827) );
  XNOR2_X1 U4012 ( .A(n3710), .B(n1530), .ZN(n1497) );
  XNOR2_X1 U4013 ( .A(n1532), .B(n1505), .ZN(n3710) );
  OAI21_X1 U4014 ( .B1(n805), .B2(n803), .A(n804), .ZN(n802) );
  INV_X1 U4015 ( .A(n803), .ZN(n1009) );
  INV_X1 U4016 ( .A(n798), .ZN(n796) );
  NAND2_X1 U4017 ( .A1(n3491), .A2(n798), .ZN(n784) );
  NOR2_X1 U4018 ( .A1(n803), .A2(n800), .ZN(n798) );
  AND2_X2 U4019 ( .A1(n3723), .A2(n3724), .ZN(n766) );
  NOR2_X1 U4020 ( .A1(n3549), .A2(n1430), .ZN(n3711) );
  NOR2_X1 U4021 ( .A1(n3698), .A2(n3097), .ZN(n3712) );
  NOR2_X1 U4022 ( .A1(n375), .A2(n3438), .ZN(n3713) );
  XNOR2_X1 U4023 ( .A(n529), .B(n327), .ZN(n3097) );
  NAND2_X1 U4024 ( .A1(n1004), .A2(n778), .ZN(n558) );
  NOR2_X1 U4025 ( .A1(n3460), .A2(n2788), .ZN(n3714) );
  NOR2_X1 U4026 ( .A1(n2787), .A2(n405), .ZN(n3715) );
  OR2_X1 U4027 ( .A1(n3714), .A2(n3715), .ZN(n2218) );
  XNOR2_X1 U4028 ( .A(n487), .B(n357), .ZN(n2788) );
  XNOR2_X1 U4029 ( .A(n489), .B(n357), .ZN(n2787) );
  NAND2_X1 U4030 ( .A1(n2547), .A2(n2323), .ZN(n3716) );
  NAND2_X1 U4031 ( .A1(n2547), .A2(n2355), .ZN(n3717) );
  NAND2_X1 U4032 ( .A1(n2323), .A2(n2355), .ZN(n3718) );
  NAND3_X1 U4033 ( .A1(n3716), .A2(n3718), .A3(n3717), .ZN(n1767) );
  OAI21_X1 U4034 ( .B1(n843), .B2(n830), .A(n3409), .ZN(n3720) );
  OR2_X1 U4035 ( .A1(n3519), .A2(n3107), .ZN(n3721) );
  OR2_X1 U4036 ( .A1(n3106), .A2(n3488), .ZN(n3722) );
  NAND2_X1 U4037 ( .A1(n3721), .A2(n3722), .ZN(n2547) );
  OAI22_X1 U4038 ( .A1(n3562), .A2(n2890), .B1(n2889), .B2(n396), .ZN(n2323)
         );
  XNOR2_X1 U4039 ( .A(n509), .B(n327), .ZN(n3107) );
  XNOR2_X1 U4040 ( .A(n511), .B(n327), .ZN(n3106) );
  NOR2_X2 U4041 ( .A1(n1918), .A2(n1933), .ZN(n887) );
  NAND2_X2 U4042 ( .A1(n1918), .A2(n1933), .ZN(n888) );
  NAND2_X2 U4043 ( .A1(n1842), .A2(n1861), .ZN(n865) );
  NOR2_X2 U4044 ( .A1(n1842), .A2(n1861), .ZN(n864) );
  NAND2_X1 U4045 ( .A1(n776), .A2(n767), .ZN(n3723) );
  INV_X1 U4046 ( .A(n768), .ZN(n3724) );
  XNOR2_X1 U4047 ( .A(n3725), .B(n2572), .ZN(n1571) );
  XNOR2_X1 U4048 ( .A(n2476), .B(n2540), .ZN(n3725) );
  BUF_X1 U4049 ( .A(n787), .Z(n3726) );
  INV_X1 U4050 ( .A(n3711), .ZN(n1003) );
  INV_X1 U4051 ( .A(n728), .ZN(n726) );
  XNOR2_X1 U4052 ( .A(n662), .B(n541), .ZN(product[54]) );
  XOR2_X1 U4053 ( .A(n2225), .B(n2577), .Z(n3727) );
  XOR2_X1 U4054 ( .A(n3727), .B(n2545), .Z(n1720) );
  XOR2_X1 U4055 ( .A(n1722), .B(n1716), .Z(n3728) );
  XOR2_X1 U4056 ( .A(n3728), .B(n1720), .Z(n1708) );
  NAND2_X1 U4057 ( .A1(n2225), .A2(n2577), .ZN(n3729) );
  NAND2_X1 U4058 ( .A1(n2225), .A2(n2545), .ZN(n3730) );
  NAND2_X1 U4059 ( .A1(n2577), .A2(n2545), .ZN(n3731) );
  NAND3_X1 U4060 ( .A1(n3729), .A2(n3730), .A3(n3731), .ZN(n1719) );
  NAND2_X1 U4061 ( .A1(n1722), .A2(n1716), .ZN(n3732) );
  NAND2_X1 U4062 ( .A1(n1722), .A2(n1720), .ZN(n3733) );
  NAND2_X1 U4063 ( .A1(n1716), .A2(n1720), .ZN(n3734) );
  NAND3_X1 U4064 ( .A1(n3732), .A2(n3733), .A3(n3734), .ZN(n1707) );
  OR2_X1 U4065 ( .A1(n3461), .A2(n2795), .ZN(n3735) );
  OR2_X1 U4066 ( .A1(n2794), .A2(n405), .ZN(n3736) );
  NAND2_X1 U4067 ( .A1(n3735), .A2(n3736), .ZN(n2225) );
  OAI21_X1 U4068 ( .B1(n811), .B2(n815), .A(n812), .ZN(n810) );
  XNOR2_X1 U4069 ( .A(n473), .B(n357), .ZN(n2795) );
  XNOR2_X1 U4070 ( .A(n475), .B(n357), .ZN(n2794) );
  OAI21_X1 U4071 ( .B1(n731), .B2(n748), .A(n732), .ZN(n730) );
  XNOR2_X1 U4072 ( .A(n771), .B(n556), .ZN(product[39]) );
  INV_X1 U4073 ( .A(n783), .ZN(n782) );
  INV_X8 U4074 ( .A(n3628), .ZN(n372) );
  NAND2_X1 U4075 ( .A1(n1545), .A2(n1543), .ZN(n3740) );
  NAND2_X1 U4076 ( .A1(n1545), .A2(n1541), .ZN(n3741) );
  NAND2_X1 U4077 ( .A1(n1543), .A2(n1541), .ZN(n3742) );
  NAND3_X2 U4078 ( .A1(n3740), .A2(n3741), .A3(n3742), .ZN(n1530) );
  NAND2_X1 U4079 ( .A1(n1532), .A2(n1505), .ZN(n3743) );
  NAND2_X1 U4080 ( .A1(n1532), .A2(n1530), .ZN(n3744) );
  NAND2_X1 U4081 ( .A1(n1505), .A2(n1530), .ZN(n3745) );
  NAND3_X1 U4082 ( .A1(n3743), .A2(n3744), .A3(n3745), .ZN(n1496) );
  XOR2_X1 U4083 ( .A(n3702), .B(n2187), .Z(n3746) );
  XOR2_X1 U4084 ( .A(n2219), .B(n3746), .Z(n1543) );
  NAND2_X1 U4085 ( .A1(n2219), .A2(n3702), .ZN(n3747) );
  NAND2_X1 U4086 ( .A1(n2219), .A2(n2187), .ZN(n3748) );
  NAND2_X1 U4087 ( .A1(n3702), .A2(n2187), .ZN(n3749) );
  NAND3_X1 U4088 ( .A1(n3747), .A2(n3749), .A3(n3748), .ZN(n1542) );
  OAI22_X1 U4089 ( .A1(n458), .A2(n2758), .B1(n2757), .B2(n3638), .ZN(n2187)
         );
  OAI22_X1 U4090 ( .A1(n3703), .A2(n3068), .B1(n3067), .B2(n3604), .ZN(n2507)
         );
  XNOR2_X1 U4091 ( .A(n650), .B(n539), .ZN(product[56]) );
  XNOR2_X1 U4092 ( .A(n643), .B(n538), .ZN(product[57]) );
  XNOR2_X1 U4093 ( .A(n698), .B(n546), .ZN(product[49]) );
  XNOR2_X1 U4094 ( .A(n595), .B(n3750), .ZN(product[63]) );
  XNOR2_X1 U4095 ( .A(n1042), .B(n1041), .ZN(n3750) );
  INV_X1 U4096 ( .A(n3496), .ZN(n685) );
  NAND2_X2 U4097 ( .A1(n1750), .A2(n1773), .ZN(n840) );
  INV_X8 U4098 ( .A(n3753), .ZN(n411) );
  AOI21_X1 U4099 ( .B1(n3665), .B2(n3663), .A(n3726), .ZN(n3756) );
  INV_X8 U4100 ( .A(n3757), .ZN(n387) );
  INV_X8 U4101 ( .A(n3759), .ZN(n399) );
  NAND2_X1 U4102 ( .A1(n1003), .A2(n3522), .ZN(n557) );
  OAI21_X1 U4103 ( .B1(n774), .B2(n3711), .A(n3522), .ZN(n771) );
  NAND2_X1 U4104 ( .A1(n1403), .A2(n1430), .ZN(n773) );
  OAI21_X1 U4105 ( .B1(n896), .B2(n883), .A(n3419), .ZN(n882) );
  INV_X1 U4106 ( .A(n3690), .ZN(n855) );
  OAI21_X1 U4107 ( .B1(n861), .B2(n865), .A(n862), .ZN(n860) );
  BUF_X1 U4108 ( .A(n775), .Z(n3765) );
  XOR2_X1 U4109 ( .A(n682), .B(n545), .Z(product[50]) );
  NAND2_X1 U4110 ( .A1(n791), .A2(n794), .ZN(n561) );
  INV_X8 U4111 ( .A(n3766), .ZN(n381) );
  OAI21_X1 U4112 ( .B1(n782), .B2(n3420), .A(n3465), .ZN(n779) );
  INV_X1 U4113 ( .A(n780), .ZN(n1005) );
  NAND2_X1 U4114 ( .A1(n3547), .A2(n817), .ZN(n807) );
  BUF_X1 U4115 ( .A(n776), .Z(n3768) );
  OAI21_X1 U4116 ( .B1(n807), .B2(n3719), .A(n808), .ZN(n3769) );
  OAI21_X2 U4117 ( .B1(n827), .B2(n807), .A(n808), .ZN(n806) );
  XOR2_X1 U4118 ( .A(n1577), .B(n1573), .Z(n3770) );
  XOR2_X1 U4119 ( .A(n3770), .B(n1571), .Z(n1563) );
  NAND2_X1 U4120 ( .A1(n2476), .A2(n2540), .ZN(n3771) );
  NAND2_X1 U4121 ( .A1(n2476), .A2(n2572), .ZN(n3772) );
  NAND2_X1 U4122 ( .A1(n2540), .A2(n2572), .ZN(n3773) );
  NAND3_X1 U4123 ( .A1(n3771), .A2(n3772), .A3(n3773), .ZN(n1570) );
  NAND2_X1 U4124 ( .A1(n1577), .A2(n1573), .ZN(n3774) );
  NAND2_X1 U4125 ( .A1(n1577), .A2(n1571), .ZN(n3775) );
  NAND2_X1 U4126 ( .A1(n1573), .A2(n1571), .ZN(n3776) );
  NAND3_X1 U4127 ( .A1(n3774), .A2(n3775), .A3(n3776), .ZN(n1562) );
  NAND2_X2 U4128 ( .A1(n832), .A2(n837), .ZN(n830) );
  BUF_X1 U4129 ( .A(n3756), .Z(n3779) );
  OAI21_X1 U4130 ( .B1(n769), .B2(n773), .A(n770), .ZN(n768) );
  NAND2_X1 U4131 ( .A1(n3464), .A2(n1402), .ZN(n770) );
  NOR2_X2 U4132 ( .A1(n1281), .A2(n1302), .ZN(n738) );
  AOI21_X2 U4133 ( .B1(n997), .B2(n3659), .A(n734), .ZN(n732) );
  NOR2_X1 U4134 ( .A1(n3519), .A2(n3100), .ZN(n3782) );
  NOR2_X1 U4135 ( .A1(n3099), .A2(n375), .ZN(n3783) );
  OR2_X1 U4136 ( .A1(n3782), .A2(n3783), .ZN(n2540) );
  XNOR2_X1 U4137 ( .A(n523), .B(n327), .ZN(n3100) );
  XNOR2_X1 U4138 ( .A(n525), .B(n327), .ZN(n3099) );
  NAND2_X2 U4139 ( .A1(n1724), .A2(n1749), .ZN(n835) );
  AOI21_X2 U4140 ( .B1(n783), .B2(n3765), .A(n3768), .ZN(n774) );
  NAND2_X1 U4141 ( .A1(n1431), .A2(n1458), .ZN(n778) );
  NAND2_X1 U4142 ( .A1(n1489), .A2(n1518), .ZN(n789) );
  XNOR2_X1 U4143 ( .A(n3578), .B(n555), .ZN(product[40]) );
  XOR2_X1 U4144 ( .A(n3550), .B(n550), .Z(product[45]) );
  AOI21_X1 U4145 ( .B1(n761), .B2(n757), .A(n758), .ZN(n756) );
  AOI21_X1 U4146 ( .B1(n761), .B2(n611), .A(n3415), .ZN(n610) );
  XNOR2_X1 U4147 ( .A(n623), .B(n536), .ZN(product[59]) );
  INV_X1 U4148 ( .A(n3553), .ZN(n797) );
  INV_X1 U4149 ( .A(n3719), .ZN(n826) );
  INV_X1 U4150 ( .A(n3709), .ZN(n1004) );
  XOR2_X1 U4151 ( .A(n3527), .B(n537), .Z(product[58]) );
  INV_X1 U4152 ( .A(n3545), .ZN(n1006) );
  NOR2_X2 U4153 ( .A1(n1459), .A2(n1488), .ZN(n780) );
  XOR2_X1 U4154 ( .A(n701), .B(n547), .Z(product[48]) );
  XNOR2_X1 U4155 ( .A(n737), .B(n551), .ZN(product[44]) );
  XOR2_X1 U4156 ( .A(n3414), .B(n552), .Z(product[43]) );
  OAI22_X1 U4157 ( .A1(n422), .A2(n3131), .B1(n3130), .B2(n372), .ZN(n2572) );
  OAI22_X1 U4158 ( .A1(n3462), .A2(n2789), .B1(n2788), .B2(n405), .ZN(n2219)
         );
  INV_X1 U4159 ( .A(n3461), .ZN(n3786) );
  OAI21_X2 U4160 ( .B1(n3618), .B2(n671), .A(n672), .ZN(n670) );
  XNOR2_X1 U4161 ( .A(n3582), .B(n548), .ZN(product[47]) );
  AOI21_X2 U4162 ( .B1(n670), .B2(n654), .A(n655), .ZN(n653) );
  XOR2_X1 U4163 ( .A(n665), .B(n542), .Z(product[53]) );
  OAI21_X1 U4164 ( .B1(n665), .B2(n663), .A(n664), .ZN(n662) );
  XNOR2_X1 U4165 ( .A(n670), .B(n543), .ZN(product[52]) );
  OAI21_X1 U4166 ( .B1(n653), .B2(n644), .A(n645), .ZN(n643) );
  OAI21_X1 U4167 ( .B1(n653), .B2(n651), .A(n652), .ZN(n650) );
  XOR2_X1 U4168 ( .A(n653), .B(n540), .Z(product[55]) );
  XNOR2_X1 U4169 ( .A(n3548), .B(n553), .ZN(product[42]) );
  XNOR2_X1 U4170 ( .A(n3694), .B(n534), .ZN(product[61]) );
  XOR2_X1 U4171 ( .A(n3508), .B(n533), .Z(product[62]) );
  INV_X2 U4172 ( .A(n594), .ZN(product[1]) );
  INV_X2 U4173 ( .A(n699), .ZN(n993) );
  INV_X2 U4174 ( .A(n696), .ZN(n992) );
  INV_X2 U4175 ( .A(n680), .ZN(n991) );
  INV_X2 U4176 ( .A(n677), .ZN(n990) );
  INV_X2 U4177 ( .A(n663), .ZN(n988) );
  INV_X2 U4178 ( .A(n660), .ZN(n987) );
  INV_X2 U4179 ( .A(n651), .ZN(n986) );
  INV_X2 U4180 ( .A(n648), .ZN(n985) );
  INV_X2 U4181 ( .A(n596), .ZN(n979) );
  INV_X2 U4182 ( .A(n978), .ZN(n976) );
  INV_X2 U4183 ( .A(n975), .ZN(n973) );
  INV_X2 U4184 ( .A(n967), .ZN(n965) );
  INV_X2 U4185 ( .A(n959), .ZN(n957) );
  INV_X2 U4186 ( .A(n955), .ZN(n954) );
  INV_X2 U4187 ( .A(n953), .ZN(n951) );
  INV_X2 U4188 ( .A(n948), .ZN(n946) );
  INV_X2 U4189 ( .A(n941), .ZN(n939) );
  INV_X2 U4190 ( .A(n937), .ZN(n936) );
  INV_X2 U4191 ( .A(n935), .ZN(n933) );
  INV_X2 U4192 ( .A(n930), .ZN(n928) );
  INV_X2 U4193 ( .A(n924), .ZN(n923) );
  INV_X2 U4194 ( .A(n915), .ZN(n914) );
  INV_X2 U4195 ( .A(n913), .ZN(n911) );
  INV_X2 U4196 ( .A(n903), .ZN(n901) );
  INV_X2 U4197 ( .A(n897), .ZN(n896) );
  INV_X2 U4198 ( .A(n891), .ZN(n893) );
  INV_X2 U4199 ( .A(n875), .ZN(n873) );
  INV_X2 U4200 ( .A(n825), .ZN(n823) );
  INV_X2 U4201 ( .A(n3769), .ZN(n805) );
  INV_X2 U4202 ( .A(n748), .ZN(n746) );
  INV_X2 U4203 ( .A(n3630), .ZN(n725) );
  INV_X2 U4204 ( .A(n719), .ZN(n721) );
  INV_X2 U4205 ( .A(n718), .ZN(n996) );
  INV_X2 U4206 ( .A(n716), .ZN(n714) );
  INV_X2 U4207 ( .A(n715), .ZN(n995) );
  INV_X2 U4208 ( .A(n712), .ZN(n710) );
  INV_X2 U4209 ( .A(n711), .ZN(n709) );
  INV_X2 U4210 ( .A(n705), .ZN(n703) );
  INV_X2 U4211 ( .A(n704), .ZN(n994) );
  INV_X2 U4212 ( .A(n691), .ZN(n689) );
  INV_X2 U4213 ( .A(n669), .ZN(n667) );
  INV_X2 U4214 ( .A(n668), .ZN(n989) );
  INV_X2 U4215 ( .A(n656), .ZN(n654) );
  INV_X2 U4216 ( .A(n647), .ZN(n645) );
  INV_X2 U4217 ( .A(n646), .ZN(n644) );
  INV_X2 U4218 ( .A(n642), .ZN(n640) );
  INV_X2 U4219 ( .A(n641), .ZN(n984) );
  INV_X2 U4220 ( .A(n633), .ZN(n631) );
  INV_X2 U4221 ( .A(n625), .ZN(n627) );
  INV_X2 U4222 ( .A(n624), .ZN(n983) );
  INV_X2 U4223 ( .A(n622), .ZN(n620) );
  INV_X2 U4224 ( .A(n621), .ZN(n982) );
  INV_X2 U4225 ( .A(n609), .ZN(n607) );
  INV_X2 U4226 ( .A(n608), .ZN(n981) );
  INV_X2 U4227 ( .A(n602), .ZN(n600) );
  INV_X2 U4228 ( .A(n601), .ZN(n980) );
  INV_X2 U4229 ( .A(n336), .ZN(n3287) );
  INV_X2 U4230 ( .A(n339), .ZN(n3286) );
  INV_X2 U4231 ( .A(n3634), .ZN(n3285) );
  INV_X2 U4232 ( .A(n3564), .ZN(n3284) );
  INV_X2 U4233 ( .A(n3645), .ZN(n3283) );
  INV_X2 U4234 ( .A(n3588), .ZN(n3282) );
  INV_X2 U4235 ( .A(n354), .ZN(n3281) );
  NAND2_X2 U4236 ( .A1(n321), .A2(n3784), .ZN(n3195) );
  NAND2_X2 U4237 ( .A1(n3778), .A2(n3784), .ZN(n3162) );
  NAND2_X2 U4238 ( .A1(n327), .A2(n3784), .ZN(n3129) );
  NAND2_X2 U4239 ( .A1(n330), .A2(n3784), .ZN(n3096) );
  NAND2_X2 U4240 ( .A1(n333), .A2(n3784), .ZN(n3063) );
  NAND2_X2 U4241 ( .A1(n336), .A2(n3784), .ZN(n3030) );
  NAND2_X2 U4242 ( .A1(n339), .A2(n3784), .ZN(n2997) );
  NAND2_X2 U4243 ( .A1(n3634), .A2(n3784), .ZN(n2964) );
  NAND2_X2 U4244 ( .A1(n3564), .A2(n3784), .ZN(n2931) );
  NAND2_X2 U4245 ( .A1(n3645), .A2(n3784), .ZN(n2898) );
  NAND2_X2 U4246 ( .A1(n3588), .A2(n3784), .ZN(n2865) );
  NAND2_X2 U4247 ( .A1(n354), .A2(n3784), .ZN(n2832) );
  NAND2_X2 U4248 ( .A1(n3467), .A2(n3784), .ZN(n2799) );
  NAND2_X2 U4249 ( .A1(n360), .A2(n3784), .ZN(n2766) );
  NAND2_X2 U4250 ( .A1(n363), .A2(n3784), .ZN(n2733) );
  NAND2_X2 U4251 ( .A1(n366), .A2(n3784), .ZN(n2700) );
  INV_X2 U4252 ( .A(n419), .ZN(n3785) );
  NOR2_X2 U4253 ( .A1(n372), .A2(n3784), .ZN(n2603) );
  NOR2_X2 U4254 ( .A1(n3488), .A2(n3784), .ZN(n2569) );
  NOR2_X2 U4255 ( .A1(n3604), .A2(n3784), .ZN(n2535) );
  NOR2_X2 U4256 ( .A1(n381), .A2(n3784), .ZN(n2501) );
  NOR2_X2 U4257 ( .A1(n3641), .A2(n3784), .ZN(n2467) );
  NOR2_X2 U4258 ( .A1(n387), .A2(n3784), .ZN(n2433) );
  NOR2_X2 U4259 ( .A1(n3650), .A2(n3784), .ZN(n2399) );
  NOR2_X2 U4260 ( .A1(n3656), .A2(n3784), .ZN(n2365) );
  NOR2_X2 U4261 ( .A1(n396), .A2(n3784), .ZN(n2331) );
  NOR2_X2 U4262 ( .A1(n399), .A2(n3784), .ZN(n2297) );
  NOR2_X2 U4263 ( .A1(n3469), .A2(n3784), .ZN(n2263) );
  NOR2_X2 U4264 ( .A1(n405), .A2(n3784), .ZN(n2229) );
  NOR2_X2 U4265 ( .A1(n3638), .A2(n3784), .ZN(n2195) );
  NOR2_X2 U4266 ( .A1(n411), .A2(n3784), .ZN(n2161) );
  INV_X2 U4267 ( .A(n1548), .ZN(n1580) );
  INV_X2 U4268 ( .A(n1486), .ZN(n1487) );
  INV_X2 U4269 ( .A(n1428), .ZN(n1429) );
  INV_X2 U4270 ( .A(n1374), .ZN(n1375) );
  INV_X2 U4271 ( .A(n1324), .ZN(n1325) );
  INV_X2 U4272 ( .A(n1278), .ZN(n1279) );
  INV_X2 U4273 ( .A(n1236), .ZN(n1237) );
  INV_X2 U4274 ( .A(n1198), .ZN(n1199) );
  INV_X2 U4275 ( .A(n1164), .ZN(n1165) );
  INV_X2 U4276 ( .A(n1134), .ZN(n1135) );
  INV_X2 U4277 ( .A(n1108), .ZN(n1109) );
  INV_X2 U4278 ( .A(n1086), .ZN(n1087) );
  INV_X2 U4279 ( .A(n1068), .ZN(n1069) );
  INV_X2 U4280 ( .A(n1054), .ZN(n1055) );
  INV_X2 U4281 ( .A(n1044), .ZN(n1045) );
  XOR2_X1 U4282 ( .A(n3787), .B(n3788), .Z(n1041) );
  XOR2_X1 U4283 ( .A(n2077), .B(n1044), .Z(n3788) );
  INV_X2 U4284 ( .A(n977), .ZN(n1040) );
  INV_X2 U4285 ( .A(n974), .ZN(n972) );
  INV_X2 U4286 ( .A(n969), .ZN(n1038) );
  INV_X2 U4287 ( .A(n966), .ZN(n964) );
  INV_X2 U4288 ( .A(n961), .ZN(n1036) );
  INV_X2 U4289 ( .A(n958), .ZN(n956) );
  INV_X2 U4290 ( .A(n952), .ZN(n950) );
  INV_X2 U4291 ( .A(n947), .ZN(n945) );
  INV_X2 U4292 ( .A(n940), .ZN(n938) );
  INV_X2 U4293 ( .A(n934), .ZN(n932) );
  INV_X2 U4294 ( .A(n929), .ZN(n927) );
  INV_X2 U4295 ( .A(n921), .ZN(n1029) );
  INV_X2 U4296 ( .A(n918), .ZN(n1028) );
  INV_X2 U4297 ( .A(n912), .ZN(n910) );
  INV_X2 U4298 ( .A(n907), .ZN(n1026) );
  INV_X2 U4299 ( .A(n902), .ZN(n900) );
  INV_X2 U4300 ( .A(n890), .ZN(n892) );
  INV_X2 U4301 ( .A(n887), .ZN(n885) );
  INV_X2 U4302 ( .A(n880), .ZN(n1022) );
  INV_X2 U4303 ( .A(n874), .ZN(n872) );
  INV_X2 U4304 ( .A(n869), .ZN(n1020) );
  INV_X2 U4305 ( .A(n861), .ZN(n1018) );
  INV_X2 U4306 ( .A(n849), .ZN(n851) );
  INV_X2 U4307 ( .A(n839), .ZN(n837) );
  INV_X2 U4308 ( .A(n834), .ZN(n832) );
  INV_X2 U4309 ( .A(n759), .ZN(n757) );
endmodule


module mul32_1_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n321, n324, n327, n330, n333, n336, n339, n342, n345, n348, n351,
         n354, n357, n360, n363, n366, n369, n372, n381, n384, n387, n390,
         n393, n396, n399, n402, n405, n408, n411, n416, n419, n422, n425,
         n428, n431, n434, n437, n443, n446, n449, n452, n455, n458, n461,
         n464, n465, n469, n471, n473, n475, n477, n479, n481, n483, n485,
         n487, n489, n491, n493, n495, n497, n499, n501, n503, n505, n507,
         n509, n511, n513, n515, n517, n519, n521, n523, n525, n527, n529,
         n531, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n600, n601, n602, n603, n604, n605, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n620, n621, n622, n623,
         n624, n625, n627, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n667, n668, n669, n670, n671, n672,
         n673, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n714, n715, n716, n717, n718, n719, n721,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n734, n735,
         n736, n737, n738, n739, n744, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n833, n835, n836, n838, n840, n841, n842, n843, n845, n847,
         n848, n849, n850, n851, n852, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1003, n1004, n1005, n1009, n1010,
         n1011, n1012, n1018, n1019, n1020, n1022, n1026, n1028, n1029, n1036,
         n1038, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3228, n3229, n3230, n3231, n3232,
         n3234, n3237, n3238, n3239, n3241, n3242, n3243, n3278, n3279, n3281,
         n3282, n3283, n3286, n3288, n3289, n3290, n3292, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755;
  assign n321 = a[1];
  assign n324 = a[3];
  assign n327 = a[5];
  assign n330 = a[7];
  assign n333 = a[9];
  assign n336 = a[11];
  assign n339 = a[13];
  assign n342 = a[15];
  assign n345 = a[17];
  assign n348 = a[19];
  assign n351 = a[21];
  assign n354 = a[23];
  assign n357 = a[25];
  assign n360 = a[27];
  assign n363 = a[29];
  assign n366 = a[31];
  assign n465 = b[0];
  assign n469 = b[1];
  assign n471 = b[2];
  assign n473 = b[3];
  assign n475 = b[4];
  assign n477 = b[5];
  assign n479 = b[6];
  assign n481 = b[7];
  assign n483 = b[8];
  assign n485 = b[9];
  assign n487 = b[10];
  assign n489 = b[11];
  assign n491 = b[12];
  assign n493 = b[13];
  assign n495 = b[14];
  assign n497 = b[15];
  assign n499 = b[16];
  assign n501 = b[17];
  assign n503 = b[18];
  assign n505 = b[19];
  assign n507 = b[20];
  assign n509 = b[21];
  assign n511 = b[22];
  assign n513 = b[23];
  assign n515 = b[24];
  assign n517 = b[25];
  assign n519 = b[26];
  assign n521 = b[27];
  assign n523 = b[28];
  assign n525 = b[29];
  assign n527 = b[30];
  assign n529 = b[31];

  NOR2_X4 U324 ( .A1(n1043), .A2(n1046), .ZN(n596) );
  NAND2_X4 U325 ( .A1(n1043), .A2(n1046), .ZN(n597) );
  NAND2_X4 U330 ( .A1(n980), .A2(n602), .ZN(n534) );
  NOR2_X4 U332 ( .A1(n1050), .A2(n1047), .ZN(n601) );
  NAND2_X4 U333 ( .A1(n1050), .A2(n1047), .ZN(n602) );
  XOR2_X2 U334 ( .A(n610), .B(n535), .Z(product[60]) );
  NAND2_X4 U340 ( .A1(n981), .A2(n609), .ZN(n535) );
  NOR2_X4 U342 ( .A1(n1051), .A2(n1056), .ZN(n608) );
  NAND2_X4 U343 ( .A1(n1051), .A2(n1056), .ZN(n609) );
  NAND2_X4 U348 ( .A1(n690), .A2(n615), .ZN(n613) );
  AOI21_X4 U349 ( .B1(n691), .B2(n615), .A(n616), .ZN(n614) );
  NOR2_X4 U350 ( .A1(n633), .A2(n617), .ZN(n615) );
  OAI21_X4 U351 ( .B1(n634), .B2(n617), .A(n618), .ZN(n616) );
  NAND2_X4 U352 ( .A1(n983), .A2(n982), .ZN(n617) );
  AOI21_X4 U353 ( .B1(n982), .B2(n627), .A(n620), .ZN(n618) );
  NAND2_X4 U356 ( .A1(n982), .A2(n622), .ZN(n536) );
  NOR2_X4 U358 ( .A1(n1057), .A2(n1062), .ZN(n621) );
  NAND2_X4 U359 ( .A1(n1057), .A2(n1062), .ZN(n622) );
  NAND2_X4 U366 ( .A1(n983), .A2(n625), .ZN(n537) );
  NOR2_X4 U368 ( .A1(n1063), .A2(n1070), .ZN(n624) );
  NAND2_X4 U369 ( .A1(n1063), .A2(n1070), .ZN(n625) );
  NAND2_X4 U374 ( .A1(n673), .A2(n635), .ZN(n633) );
  AOI21_X4 U375 ( .B1(n635), .B2(n676), .A(n636), .ZN(n634) );
  NOR2_X4 U376 ( .A1(n656), .A2(n637), .ZN(n635) );
  NAND2_X4 U378 ( .A1(n646), .A2(n984), .ZN(n637) );
  AOI21_X4 U379 ( .B1(n647), .B2(n984), .A(n640), .ZN(n638) );
  NAND2_X4 U382 ( .A1(n984), .A2(n642), .ZN(n538) );
  NOR2_X4 U384 ( .A1(n1071), .A2(n1078), .ZN(n641) );
  NAND2_X4 U385 ( .A1(n1071), .A2(n1078), .ZN(n642) );
  NOR2_X4 U390 ( .A1(n651), .A2(n648), .ZN(n646) );
  OAI21_X4 U391 ( .B1(n648), .B2(n652), .A(n649), .ZN(n647) );
  NAND2_X4 U392 ( .A1(n985), .A2(n649), .ZN(n539) );
  NOR2_X4 U394 ( .A1(n1079), .A2(n1088), .ZN(n648) );
  NAND2_X4 U395 ( .A1(n1079), .A2(n1088), .ZN(n649) );
  NAND2_X4 U398 ( .A1(n986), .A2(n652), .ZN(n540) );
  NOR2_X4 U400 ( .A1(n1089), .A2(n1098), .ZN(n651) );
  NAND2_X4 U401 ( .A1(n1089), .A2(n1098), .ZN(n652) );
  NAND2_X4 U406 ( .A1(n658), .A2(n989), .ZN(n656) );
  AOI21_X4 U407 ( .B1(n658), .B2(n667), .A(n659), .ZN(n657) );
  NOR2_X4 U408 ( .A1(n663), .A2(n660), .ZN(n658) );
  OAI21_X4 U409 ( .B1(n660), .B2(n664), .A(n661), .ZN(n659) );
  NAND2_X4 U410 ( .A1(n987), .A2(n661), .ZN(n541) );
  NOR2_X4 U412 ( .A1(n1099), .A2(n1110), .ZN(n660) );
  NAND2_X4 U413 ( .A1(n1099), .A2(n1110), .ZN(n661) );
  NAND2_X4 U416 ( .A1(n988), .A2(n664), .ZN(n542) );
  NOR2_X4 U418 ( .A1(n1111), .A2(n1122), .ZN(n663) );
  NAND2_X4 U419 ( .A1(n1111), .A2(n1122), .ZN(n664) );
  NAND2_X4 U424 ( .A1(n989), .A2(n669), .ZN(n543) );
  XNOR2_X2 U428 ( .A(n679), .B(n544), .ZN(product[51]) );
  NAND2_X4 U430 ( .A1(n686), .A2(n673), .ZN(n671) );
  NOR2_X4 U434 ( .A1(n680), .A2(n677), .ZN(n673) );
  NAND2_X4 U436 ( .A1(n990), .A2(n678), .ZN(n544) );
  NOR2_X4 U438 ( .A1(n1137), .A2(n1150), .ZN(n677) );
  NAND2_X4 U439 ( .A1(n1137), .A2(n1150), .ZN(n678) );
  XOR2_X2 U440 ( .A(n682), .B(n545), .Z(product[50]) );
  OAI21_X4 U441 ( .B1(n682), .B2(n680), .A(n681), .ZN(n679) );
  NAND2_X4 U442 ( .A1(n991), .A2(n681), .ZN(n545) );
  NOR2_X4 U444 ( .A1(n1151), .A2(n1166), .ZN(n680) );
  NAND2_X4 U445 ( .A1(n1151), .A2(n1166), .ZN(n681) );
  NOR2_X4 U451 ( .A1(n727), .A2(n688), .ZN(n686) );
  NOR2_X4 U455 ( .A1(n692), .A2(n711), .ZN(n690) );
  OAI21_X4 U456 ( .B1(n692), .B2(n712), .A(n693), .ZN(n691) );
  NOR2_X4 U459 ( .A1(n699), .A2(n696), .ZN(n694) );
  NAND2_X4 U461 ( .A1(n992), .A2(n697), .ZN(n546) );
  NOR2_X4 U463 ( .A1(n1167), .A2(n1182), .ZN(n696) );
  NAND2_X4 U467 ( .A1(n993), .A2(n700), .ZN(n547) );
  NOR2_X4 U469 ( .A1(n1183), .A2(n1200), .ZN(n699) );
  NAND2_X4 U470 ( .A1(n1183), .A2(n1200), .ZN(n700) );
  NAND2_X4 U475 ( .A1(n994), .A2(n705), .ZN(n548) );
  NOR2_X4 U477 ( .A1(n1201), .A2(n1218), .ZN(n704) );
  NAND2_X4 U478 ( .A1(n1201), .A2(n1218), .ZN(n705) );
  NAND2_X4 U481 ( .A1(n725), .A2(n709), .ZN(n707) );
  AOI21_X4 U486 ( .B1(n995), .B2(n721), .A(n714), .ZN(n712) );
  NAND2_X4 U489 ( .A1(n995), .A2(n716), .ZN(n549) );
  NAND2_X4 U499 ( .A1(n996), .A2(n719), .ZN(n550) );
  NOR2_X4 U501 ( .A1(n1239), .A2(n1258), .ZN(n718) );
  NAND2_X4 U502 ( .A1(n1239), .A2(n1258), .ZN(n719) );
  NAND2_X4 U533 ( .A1(n999), .A2(n748), .ZN(n553) );
  XOR2_X2 U537 ( .A(n756), .B(n554), .Z(product[41]) );
  NAND2_X4 U543 ( .A1(n3447), .A2(n755), .ZN(n554) );
  XNOR2_X2 U555 ( .A(n771), .B(n556), .ZN(product[39]) );
  XOR2_X2 U588 ( .A(n790), .B(n560), .Z(product[35]) );
  NAND2_X4 U595 ( .A1(n3701), .A2(n789), .ZN(n560) );
  XNOR2_X2 U599 ( .A(n795), .B(n561), .ZN(product[34]) );
  AOI21_X4 U600 ( .B1(n795), .B2(n791), .A(n792), .ZN(n790) );
  XNOR2_X2 U607 ( .A(n802), .B(n562), .ZN(product[33]) );
  XNOR2_X2 U623 ( .A(n813), .B(n564), .ZN(product[31]) );
  XOR2_X2 U634 ( .A(n816), .B(n565), .Z(product[30]) );
  XOR2_X2 U640 ( .A(n821), .B(n566), .Z(product[29]) );
  NAND2_X4 U644 ( .A1(n1012), .A2(n820), .ZN(n566) );
  XNOR2_X2 U648 ( .A(n826), .B(n567), .ZN(product[28]) );
  AOI21_X4 U649 ( .B1(n826), .B2(n822), .A(n823), .ZN(n821) );
  NAND2_X4 U652 ( .A1(n822), .A2(n825), .ZN(n567) );
  XOR2_X2 U656 ( .A(n836), .B(n568), .Z(product[27]) );
  NAND2_X4 U665 ( .A1(n3665), .A2(n835), .ZN(n568) );
  XNOR2_X2 U669 ( .A(n841), .B(n569), .ZN(product[26]) );
  AOI21_X4 U670 ( .B1(n841), .B2(n3679), .A(n838), .ZN(n836) );
  XNOR2_X2 U677 ( .A(n848), .B(n570), .ZN(product[25]) );
  XOR2_X2 U687 ( .A(n855), .B(n571), .Z(product[24]) );
  XNOR2_X2 U697 ( .A(n863), .B(n572), .ZN(product[23]) );
  NAND2_X4 U704 ( .A1(n1018), .A2(n862), .ZN(n572) );
  XOR2_X2 U708 ( .A(n866), .B(n573), .Z(product[22]) );
  NAND2_X4 U710 ( .A1(n1019), .A2(n865), .ZN(n573) );
  XOR2_X2 U714 ( .A(n871), .B(n574), .Z(product[21]) );
  OAI21_X4 U717 ( .B1(n869), .B2(n875), .A(n870), .ZN(n868) );
  NAND2_X4 U718 ( .A1(n1020), .A2(n870), .ZN(n574) );
  XNOR2_X2 U722 ( .A(n876), .B(n575), .ZN(product[20]) );
  AOI21_X4 U723 ( .B1(n876), .B2(n872), .A(n873), .ZN(n871) );
  NAND2_X4 U726 ( .A1(n872), .A2(n875), .ZN(n575) );
  NAND2_X4 U729 ( .A1(n1882), .A2(n1899), .ZN(n875) );
  XNOR2_X2 U730 ( .A(n882), .B(n576), .ZN(product[19]) );
  NAND2_X4 U735 ( .A1(n1022), .A2(n881), .ZN(n576) );
  NOR2_X4 U737 ( .A1(n1900), .A2(n1917), .ZN(n880) );
  NAND2_X4 U738 ( .A1(n1900), .A2(n1917), .ZN(n881) );
  XNOR2_X2 U739 ( .A(n889), .B(n577), .ZN(product[18]) );
  XOR2_X2 U749 ( .A(n896), .B(n578), .Z(product[17]) );
  OAI21_X4 U750 ( .B1(n896), .B2(n890), .A(n891), .ZN(n889) );
  NAND2_X4 U755 ( .A1(n892), .A2(n891), .ZN(n578) );
  XOR2_X2 U759 ( .A(n904), .B(n579), .Z(product[16]) );
  NAND2_X4 U766 ( .A1(n900), .A2(n903), .ZN(n579) );
  NOR2_X4 U768 ( .A1(n1950), .A2(n1963), .ZN(n902) );
  NAND2_X4 U769 ( .A1(n1950), .A2(n1963), .ZN(n903) );
  XOR2_X2 U770 ( .A(n909), .B(n580), .Z(product[15]) );
  AOI21_X4 U771 ( .B1(n914), .B2(n905), .A(n906), .ZN(n904) );
  NOR2_X4 U772 ( .A1(n907), .A2(n912), .ZN(n905) );
  NAND2_X4 U774 ( .A1(n1026), .A2(n908), .ZN(n580) );
  NOR2_X4 U776 ( .A1(n1964), .A2(n1977), .ZN(n907) );
  XNOR2_X2 U778 ( .A(n914), .B(n581), .ZN(product[14]) );
  AOI21_X4 U779 ( .B1(n914), .B2(n910), .A(n911), .ZN(n909) );
  NAND2_X4 U782 ( .A1(n910), .A2(n913), .ZN(n581) );
  NOR2_X4 U784 ( .A1(n1978), .A2(n1989), .ZN(n912) );
  NAND2_X4 U785 ( .A1(n1978), .A2(n1989), .ZN(n913) );
  XNOR2_X2 U786 ( .A(n920), .B(n582), .ZN(product[13]) );
  AOI21_X4 U788 ( .B1(n916), .B2(n924), .A(n917), .ZN(n915) );
  NOR2_X4 U789 ( .A1(n918), .A2(n921), .ZN(n916) );
  OAI21_X4 U790 ( .B1(n918), .B2(n922), .A(n919), .ZN(n917) );
  NAND2_X4 U791 ( .A1(n1028), .A2(n919), .ZN(n582) );
  NOR2_X4 U793 ( .A1(n1990), .A2(n2001), .ZN(n918) );
  NAND2_X4 U794 ( .A1(n1990), .A2(n2001), .ZN(n919) );
  XOR2_X2 U795 ( .A(n923), .B(n583), .Z(product[12]) );
  OAI21_X4 U796 ( .B1(n923), .B2(n921), .A(n922), .ZN(n920) );
  NAND2_X4 U797 ( .A1(n1029), .A2(n922), .ZN(n583) );
  NOR2_X4 U799 ( .A1(n2002), .A2(n2011), .ZN(n921) );
  NAND2_X4 U800 ( .A1(n2002), .A2(n2011), .ZN(n922) );
  XOR2_X2 U801 ( .A(n931), .B(n584), .Z(product[11]) );
  OAI21_X4 U803 ( .B1(n925), .B2(n937), .A(n926), .ZN(n924) );
  NAND2_X4 U804 ( .A1(n932), .A2(n927), .ZN(n925) );
  AOI21_X4 U805 ( .B1(n927), .B2(n933), .A(n928), .ZN(n926) );
  NAND2_X4 U808 ( .A1(n927), .A2(n930), .ZN(n584) );
  NOR2_X4 U810 ( .A1(n2012), .A2(n2021), .ZN(n929) );
  NAND2_X4 U811 ( .A1(n2012), .A2(n2021), .ZN(n930) );
  XNOR2_X2 U812 ( .A(n585), .B(n936), .ZN(product[10]) );
  AOI21_X4 U813 ( .B1(n936), .B2(n932), .A(n933), .ZN(n931) );
  NAND2_X4 U816 ( .A1(n932), .A2(n935), .ZN(n585) );
  NOR2_X4 U818 ( .A1(n2022), .A2(n2029), .ZN(n934) );
  NAND2_X4 U819 ( .A1(n2022), .A2(n2029), .ZN(n935) );
  XNOR2_X2 U820 ( .A(n586), .B(n942), .ZN(product[9]) );
  AOI21_X4 U822 ( .B1(n942), .B2(n938), .A(n939), .ZN(n937) );
  NAND2_X4 U825 ( .A1(n938), .A2(n941), .ZN(n586) );
  NOR2_X4 U827 ( .A1(n2030), .A2(n2037), .ZN(n940) );
  NAND2_X4 U828 ( .A1(n2030), .A2(n2037), .ZN(n941) );
  XOR2_X2 U829 ( .A(n949), .B(n587), .Z(product[8]) );
  OAI21_X4 U830 ( .B1(n943), .B2(n955), .A(n944), .ZN(n942) );
  NAND2_X4 U831 ( .A1(n945), .A2(n950), .ZN(n943) );
  AOI21_X4 U832 ( .B1(n945), .B2(n951), .A(n946), .ZN(n944) );
  NAND2_X4 U835 ( .A1(n945), .A2(n948), .ZN(n587) );
  NOR2_X4 U837 ( .A1(n2038), .A2(n2043), .ZN(n947) );
  NAND2_X4 U838 ( .A1(n2038), .A2(n2043), .ZN(n948) );
  XNOR2_X2 U839 ( .A(n954), .B(n588), .ZN(product[7]) );
  AOI21_X4 U840 ( .B1(n954), .B2(n950), .A(n951), .ZN(n949) );
  NAND2_X4 U843 ( .A1(n950), .A2(n953), .ZN(n588) );
  NOR2_X4 U845 ( .A1(n2044), .A2(n2049), .ZN(n952) );
  NAND2_X4 U846 ( .A1(n2044), .A2(n2049), .ZN(n953) );
  XNOR2_X2 U847 ( .A(n589), .B(n960), .ZN(product[6]) );
  AOI21_X4 U849 ( .B1(n956), .B2(n960), .A(n957), .ZN(n955) );
  NAND2_X4 U852 ( .A1(n956), .A2(n959), .ZN(n589) );
  NOR2_X4 U854 ( .A1(n2050), .A2(n2053), .ZN(n958) );
  NAND2_X4 U855 ( .A1(n2050), .A2(n2053), .ZN(n959) );
  XOR2_X2 U856 ( .A(n590), .B(n963), .Z(product[5]) );
  OAI21_X4 U857 ( .B1(n961), .B2(n963), .A(n962), .ZN(n960) );
  NAND2_X4 U858 ( .A1(n1036), .A2(n962), .ZN(n590) );
  NOR2_X4 U860 ( .A1(n2054), .A2(n2057), .ZN(n961) );
  NAND2_X4 U861 ( .A1(n2054), .A2(n2057), .ZN(n962) );
  XNOR2_X2 U862 ( .A(n591), .B(n968), .ZN(product[4]) );
  AOI21_X4 U863 ( .B1(n964), .B2(n968), .A(n965), .ZN(n963) );
  NAND2_X4 U866 ( .A1(n964), .A2(n967), .ZN(n591) );
  NOR2_X4 U868 ( .A1(n2058), .A2(n2059), .ZN(n966) );
  NAND2_X4 U869 ( .A1(n2058), .A2(n2059), .ZN(n967) );
  XOR2_X2 U870 ( .A(n592), .B(n971), .Z(product[3]) );
  OAI21_X4 U871 ( .B1(n969), .B2(n971), .A(n970), .ZN(n968) );
  NAND2_X4 U872 ( .A1(n1038), .A2(n970), .ZN(n592) );
  NOR2_X4 U874 ( .A1(n2060), .A2(n2075), .ZN(n969) );
  NAND2_X4 U875 ( .A1(n2060), .A2(n2075), .ZN(n970) );
  XNOR2_X2 U876 ( .A(n593), .B(n976), .ZN(product[2]) );
  AOI21_X4 U877 ( .B1(n972), .B2(n976), .A(n973), .ZN(n971) );
  NAND2_X4 U880 ( .A1(n972), .A2(n975), .ZN(n593) );
  NOR2_X4 U882 ( .A1(n2603), .A2(n2635), .ZN(n974) );
  NAND2_X4 U883 ( .A1(n2603), .A2(n2635), .ZN(n975) );
  NAND2_X4 U886 ( .A1(n1040), .A2(n978), .ZN(n594) );
  NOR2_X4 U888 ( .A1(n2636), .A2(n2076), .ZN(n977) );
  NAND2_X4 U889 ( .A1(n2636), .A2(n2076), .ZN(n978) );
  FA_X1 U890 ( .A(n2095), .B(n1045), .CI(n1048), .CO(n1042), .S(n1043) );
  FA_X1 U892 ( .A(n1052), .B(n2128), .CI(n1049), .CO(n1046), .S(n1047) );
  FA_X1 U893 ( .A(n2078), .B(n1054), .CI(n2096), .CO(n1048), .S(n1049) );
  FA_X1 U894 ( .A(n1053), .B(n1060), .CI(n1058), .CO(n1050), .S(n1051) );
  FA_X1 U895 ( .A(n2129), .B(n1055), .CI(n2097), .CO(n1052), .S(n1053) );
  FA_X1 U897 ( .A(n1064), .B(n1061), .CI(n1059), .CO(n1056), .S(n1057) );
  FA_X1 U898 ( .A(n2162), .B(n2098), .CI(n1066), .CO(n1058), .S(n1059) );
  FA_X1 U899 ( .A(n2079), .B(n1068), .CI(n2130), .CO(n1060), .S(n1061) );
  FA_X1 U900 ( .A(n1072), .B(n1067), .CI(n1065), .CO(n1062), .S(n1063) );
  FA_X1 U901 ( .A(n1076), .B(n2099), .CI(n1074), .CO(n1064), .S(n1065) );
  FA_X1 U902 ( .A(n2163), .B(n1069), .CI(n2131), .CO(n1066), .S(n1067) );
  FA_X1 U904 ( .A(n1080), .B(n1082), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U905 ( .A(n1077), .B(n1084), .CI(n1075), .CO(n1072), .S(n1073) );
  FA_X1 U906 ( .A(n2132), .B(n2100), .CI(n2196), .CO(n1074), .S(n1075) );
  FA_X1 U907 ( .A(n2080), .B(n1086), .CI(n2164), .CO(n1076), .S(n1077) );
  FA_X1 U908 ( .A(n1090), .B(n1083), .CI(n1081), .CO(n1078), .S(n1079) );
  FA_X1 U909 ( .A(n1085), .B(n1094), .CI(n1092), .CO(n1080), .S(n1081) );
  FA_X1 U910 ( .A(n2101), .B(n2133), .CI(n1096), .CO(n1082), .S(n1083) );
  FA_X1 U911 ( .A(n2197), .B(n1087), .CI(n2165), .CO(n1084), .S(n1085) );
  FA_X1 U913 ( .A(n1100), .B(n1093), .CI(n1091), .CO(n1088), .S(n1089) );
  FA_X1 U914 ( .A(n1095), .B(n1097), .CI(n1102), .CO(n1090), .S(n1091) );
  FA_X1 U915 ( .A(n1106), .B(n2230), .CI(n1104), .CO(n1092), .S(n1093) );
  FA_X1 U916 ( .A(n2102), .B(n2134), .CI(n2198), .CO(n1094), .S(n1095) );
  FA_X1 U917 ( .A(n2081), .B(n1108), .CI(n2166), .CO(n1096), .S(n1097) );
  FA_X1 U918 ( .A(n1112), .B(n1103), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U919 ( .A(n1116), .B(n1105), .CI(n1114), .CO(n1100), .S(n1101) );
  FA_X1 U920 ( .A(n1118), .B(n1120), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U921 ( .A(n2135), .B(n2103), .CI(n2167), .CO(n1104), .S(n1105) );
  FA_X1 U922 ( .A(n2231), .B(n1109), .CI(n2199), .CO(n1106), .S(n1107) );
  FA_X1 U924 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U925 ( .A(n1117), .B(n1128), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U926 ( .A(n1121), .B(n1130), .CI(n1119), .CO(n1114), .S(n1115) );
  FA_X1 U927 ( .A(n2264), .B(n2136), .CI(n1132), .CO(n1116), .S(n1117) );
  FA_X1 U928 ( .A(n2104), .B(n2168), .CI(n2232), .CO(n1118), .S(n1119) );
  FA_X1 U929 ( .A(n2082), .B(n1134), .CI(n2200), .CO(n1120), .S(n1121) );
  FA_X1 U930 ( .A(n1138), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U931 ( .A(n1129), .B(n1142), .CI(n1140), .CO(n1124), .S(n1125) );
  FA_X1 U932 ( .A(n1133), .B(n1144), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U933 ( .A(n1148), .B(n2137), .CI(n1146), .CO(n1128), .S(n1129) );
  FA_X1 U934 ( .A(n2105), .B(n2201), .CI(n2169), .CO(n1130), .S(n1131) );
  FA_X1 U935 ( .A(n2265), .B(n1135), .CI(n2233), .CO(n1132), .S(n1133) );
  FA_X1 U937 ( .A(n1152), .B(n1141), .CI(n1139), .CO(n1136), .S(n1137) );
  FA_X1 U938 ( .A(n1143), .B(n1156), .CI(n1154), .CO(n1138), .S(n1139) );
  FA_X1 U939 ( .A(n1145), .B(n1147), .CI(n1158), .CO(n1140), .S(n1141) );
  FA_X1 U940 ( .A(n1160), .B(n1162), .CI(n1149), .CO(n1142), .S(n1143) );
  FA_X1 U941 ( .A(n2266), .B(n2106), .CI(n2298), .CO(n1144), .S(n1145) );
  FA_X1 U942 ( .A(n2138), .B(n2170), .CI(n2234), .CO(n1146), .S(n1147) );
  FA_X1 U943 ( .A(n2083), .B(n1164), .CI(n2202), .CO(n1148), .S(n1149) );
  FA_X1 U944 ( .A(n1168), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U945 ( .A(n1157), .B(n1172), .CI(n1170), .CO(n1152), .S(n1153) );
  FA_X1 U946 ( .A(n1174), .B(n1161), .CI(n1159), .CO(n1154), .S(n1155) );
  FA_X1 U947 ( .A(n1176), .B(n1178), .CI(n1163), .CO(n1156), .S(n1157) );
  FA_X1 U948 ( .A(n2171), .B(n2203), .CI(n1180), .CO(n1158), .S(n1159) );
  FA_X1 U949 ( .A(n2107), .B(n2235), .CI(n2139), .CO(n1160), .S(n1161) );
  FA_X1 U950 ( .A(n2299), .B(n1165), .CI(n2267), .CO(n1162), .S(n1163) );
  FA_X1 U952 ( .A(n1184), .B(n1171), .CI(n1169), .CO(n1166), .S(n1167) );
  FA_X1 U953 ( .A(n1173), .B(n1188), .CI(n1186), .CO(n1168), .S(n1169) );
  FA_X1 U954 ( .A(n1190), .B(n1179), .CI(n1175), .CO(n1170), .S(n1171) );
  FA_X1 U955 ( .A(n1181), .B(n1192), .CI(n1177), .CO(n1172), .S(n1173) );
  FA_X1 U956 ( .A(n1196), .B(n2332), .CI(n1194), .CO(n1174), .S(n1175) );
  FA_X1 U957 ( .A(n2268), .B(n2140), .CI(n2300), .CO(n1176), .S(n1177) );
  FA_X1 U958 ( .A(n2108), .B(n2204), .CI(n2172), .CO(n1178), .S(n1179) );
  FA_X1 U959 ( .A(n2084), .B(n1198), .CI(n2236), .CO(n1180), .S(n1181) );
  FA_X1 U960 ( .A(n1202), .B(n1187), .CI(n1185), .CO(n1182), .S(n1183) );
  FA_X1 U961 ( .A(n1189), .B(n1206), .CI(n1204), .CO(n1184), .S(n1185) );
  FA_X1 U962 ( .A(n1208), .B(n1210), .CI(n1191), .CO(n1186), .S(n1187) );
  FA_X1 U963 ( .A(n1193), .B(n1197), .CI(n1195), .CO(n1188), .S(n1189) );
  FA_X1 U964 ( .A(n1214), .B(n1216), .CI(n1212), .CO(n1190), .S(n1191) );
  FA_X1 U965 ( .A(n2141), .B(n2205), .CI(n2173), .CO(n1192), .S(n1193) );
  FA_X1 U966 ( .A(n2109), .B(n2269), .CI(n2237), .CO(n1194), .S(n1195) );
  FA_X1 U967 ( .A(n2333), .B(n1199), .CI(n2301), .CO(n1196), .S(n1197) );
  FA_X1 U969 ( .A(n1220), .B(n1205), .CI(n1203), .CO(n1200), .S(n1201) );
  FA_X1 U970 ( .A(n1207), .B(n1224), .CI(n1222), .CO(n1202), .S(n1203) );
  FA_X1 U971 ( .A(n1211), .B(n1226), .CI(n1209), .CO(n1204), .S(n1205) );
  FA_X1 U972 ( .A(n1215), .B(n1213), .CI(n1228), .CO(n1206), .S(n1207) );
  FA_X1 U973 ( .A(n1230), .B(n1232), .CI(n1217), .CO(n1208), .S(n1209) );
  FA_X1 U974 ( .A(n2366), .B(n2334), .CI(n1234), .CO(n1210), .S(n1211) );
  FA_X1 U975 ( .A(n2302), .B(n2174), .CI(n2270), .CO(n1212), .S(n1213) );
  FA_X1 U976 ( .A(n2142), .B(n2206), .CI(n2110), .CO(n1214), .S(n1215) );
  FA_X1 U977 ( .A(n2085), .B(n1236), .CI(n2238), .CO(n1216), .S(n1217) );
  FA_X1 U978 ( .A(n1240), .B(n1223), .CI(n1221), .CO(n1218), .S(n1219) );
  FA_X1 U979 ( .A(n1225), .B(n1244), .CI(n1242), .CO(n1220), .S(n1221) );
  FA_X1 U980 ( .A(n1246), .B(n1229), .CI(n1227), .CO(n1222), .S(n1223) );
  FA_X1 U981 ( .A(n1233), .B(n1231), .CI(n1248), .CO(n1224), .S(n1225) );
  FA_X1 U982 ( .A(n1250), .B(n1252), .CI(n1235), .CO(n1226), .S(n1227) );
  FA_X1 U983 ( .A(n1256), .B(n2239), .CI(n1254), .CO(n1228), .S(n1229) );
  FA_X1 U984 ( .A(n2175), .B(n2271), .CI(n2207), .CO(n1230), .S(n1231) );
  FA_X1 U985 ( .A(n2111), .B(n2303), .CI(n2143), .CO(n1232), .S(n1233) );
  FA_X1 U986 ( .A(n2367), .B(n1237), .CI(n2335), .CO(n1234), .S(n1235) );
  FA_X1 U988 ( .A(n1260), .B(n1243), .CI(n1241), .CO(n1238), .S(n1239) );
  FA_X1 U989 ( .A(n1245), .B(n1264), .CI(n1262), .CO(n1240), .S(n1241) );
  FA_X1 U990 ( .A(n1249), .B(n1266), .CI(n1247), .CO(n1242), .S(n1243) );
  FA_X1 U991 ( .A(n1270), .B(n1251), .CI(n1268), .CO(n1244), .S(n1245) );
  FA_X1 U992 ( .A(n1253), .B(n1257), .CI(n1255), .CO(n1246), .S(n1247) );
  FA_X1 U993 ( .A(n1272), .B(n1276), .CI(n1274), .CO(n1248), .S(n1249) );
  FA_X1 U994 ( .A(n2336), .B(n2368), .CI(n2400), .CO(n1250), .S(n1251) );
  FA_X1 U995 ( .A(n2304), .B(n2144), .CI(n2208), .CO(n1252), .S(n1253) );
  FA_X1 U996 ( .A(n2112), .B(n2240), .CI(n2176), .CO(n1254), .S(n1255) );
  FA_X1 U997 ( .A(n2086), .B(n1278), .CI(n2272), .CO(n1256), .S(n1257) );
  FA_X1 U998 ( .A(n1263), .B(n1282), .CI(n1261), .CO(n1258), .S(n1259) );
  FA_X1 U999 ( .A(n1265), .B(n1286), .CI(n1284), .CO(n1260), .S(n1261) );
  FA_X1 U1000 ( .A(n1269), .B(n1288), .CI(n1267), .CO(n1262), .S(n1263) );
  FA_X1 U1001 ( .A(n1271), .B(n1292), .CI(n1290), .CO(n1264), .S(n1265) );
  FA_X1 U1002 ( .A(n1273), .B(n1277), .CI(n1275), .CO(n1266), .S(n1267) );
  FA_X1 U1003 ( .A(n1294), .B(n1298), .CI(n1296), .CO(n1268), .S(n1269) );
  FA_X1 U1004 ( .A(n2273), .B(n2305), .CI(n1300), .CO(n1270), .S(n1271) );
  FA_X1 U1005 ( .A(n2177), .B(n2241), .CI(n2209), .CO(n1272), .S(n1273) );
  FA_X1 U1006 ( .A(n2113), .B(n2337), .CI(n2145), .CO(n1274), .S(n1275) );
  FA_X1 U1007 ( .A(n2401), .B(n1279), .CI(n2369), .CO(n1276), .S(n1277) );
  FA_X1 U1010 ( .A(n1287), .B(n1308), .CI(n1306), .CO(n1282), .S(n1283) );
  FA_X1 U1011 ( .A(n1310), .B(n1291), .CI(n1289), .CO(n1284), .S(n1285) );
  FA_X1 U1012 ( .A(n1312), .B(n1314), .CI(n1293), .CO(n1286), .S(n1287) );
  FA_X1 U1013 ( .A(n1299), .B(n1295), .CI(n1297), .CO(n1288), .S(n1289) );
  FA_X1 U1014 ( .A(n1316), .B(n1318), .CI(n1301), .CO(n1290), .S(n1291) );
  FA_X1 U1015 ( .A(n1322), .B(n2434), .CI(n1320), .CO(n1292), .S(n1293) );
  FA_X1 U1016 ( .A(n2210), .B(n2402), .CI(n2370), .CO(n1294), .S(n1295) );
  FA_X1 U1017 ( .A(n2178), .B(n2306), .CI(n2338), .CO(n1296), .S(n1297) );
  FA_X1 U1018 ( .A(n2114), .B(n2242), .CI(n2146), .CO(n1298), .S(n1299) );
  FA_X1 U1019 ( .A(n2087), .B(n1324), .CI(n2274), .CO(n1300), .S(n1301) );
  FA_X1 U1020 ( .A(n1328), .B(n1307), .CI(n1305), .CO(n1302), .S(n1303) );
  FA_X1 U1021 ( .A(n1309), .B(n1332), .CI(n1330), .CO(n1304), .S(n1305) );
  FA_X1 U1022 ( .A(n1334), .B(n1313), .CI(n1311), .CO(n1306), .S(n1307) );
  FA_X1 U1023 ( .A(n1315), .B(n1338), .CI(n1336), .CO(n1308), .S(n1309) );
  FA_X1 U1024 ( .A(n1321), .B(n1319), .CI(n1340), .CO(n1310), .S(n1311) );
  FA_X1 U1025 ( .A(n1323), .B(n1342), .CI(n1317), .CO(n1312), .S(n1313) );
  FA_X1 U1026 ( .A(n1346), .B(n1348), .CI(n1344), .CO(n1314), .S(n1315) );
  FA_X1 U1027 ( .A(n2243), .B(n2307), .CI(n2275), .CO(n1316), .S(n1317) );
  FA_X1 U1028 ( .A(n2339), .B(n2179), .CI(n2211), .CO(n1318), .S(n1319) );
  FA_X1 U1029 ( .A(n2115), .B(n2371), .CI(n2147), .CO(n1320), .S(n1321) );
  FA_X1 U1030 ( .A(n2435), .B(n1325), .CI(n2403), .CO(n1322), .S(n1323) );
  FA_X1 U1032 ( .A(n1352), .B(n1331), .CI(n1329), .CO(n1326), .S(n1327) );
  FA_X1 U1033 ( .A(n1333), .B(n1356), .CI(n1354), .CO(n1328), .S(n1329) );
  FA_X1 U1034 ( .A(n1358), .B(n1337), .CI(n1335), .CO(n1330), .S(n1331) );
  FA_X1 U1035 ( .A(n1360), .B(n1341), .CI(n1339), .CO(n1332), .S(n1333) );
  FA_X1 U1036 ( .A(n1364), .B(n1347), .CI(n1362), .CO(n1334), .S(n1335) );
  FA_X1 U1037 ( .A(n1343), .B(n1349), .CI(n1345), .CO(n1336), .S(n1337) );
  FA_X1 U1038 ( .A(n1366), .B(n1370), .CI(n1368), .CO(n1338), .S(n1339) );
  FA_X1 U1039 ( .A(n2468), .B(n2436), .CI(n1372), .CO(n1340), .S(n1341) );
  FA_X1 U1040 ( .A(n2212), .B(n2404), .CI(n2372), .CO(n1342), .S(n1343) );
  FA_X1 U1041 ( .A(n2116), .B(n2340), .CI(n2244), .CO(n1344), .S(n1345) );
  FA_X1 U1042 ( .A(n2148), .B(n2276), .CI(n2180), .CO(n1346), .S(n1347) );
  FA_X1 U1043 ( .A(n2088), .B(n1374), .CI(n2308), .CO(n1348), .S(n1349) );
  FA_X1 U1044 ( .A(n1378), .B(n1355), .CI(n1353), .CO(n1350), .S(n1351) );
  FA_X1 U1045 ( .A(n1357), .B(n1382), .CI(n1380), .CO(n1352), .S(n1353) );
  FA_X1 U1046 ( .A(n1384), .B(n1361), .CI(n1359), .CO(n1354), .S(n1355) );
  FA_X1 U1047 ( .A(n1386), .B(n1365), .CI(n1363), .CO(n1356), .S(n1357) );
  FA_X1 U1048 ( .A(n1390), .B(n1369), .CI(n1388), .CO(n1358), .S(n1359) );
  FA_X1 U1049 ( .A(n1367), .B(n1373), .CI(n1371), .CO(n1360), .S(n1361) );
  FA_X1 U1050 ( .A(n1394), .B(n1396), .CI(n1392), .CO(n1362), .S(n1363) );
  FA_X1 U1051 ( .A(n1400), .B(n2341), .CI(n1398), .CO(n1364), .S(n1365) );
  FA_X1 U1052 ( .A(n2245), .B(n2373), .CI(n2309), .CO(n1366), .S(n1367) );
  FA_X1 U1053 ( .A(n2181), .B(n2405), .CI(n2213), .CO(n1368), .S(n1369) );
  FA_X1 U1054 ( .A(n2117), .B(n2437), .CI(n2149), .CO(n1370), .S(n1371) );
  FA_X1 U1055 ( .A(n2277), .B(n1375), .CI(n2469), .CO(n1372), .S(n1373) );
  FA_X1 U1057 ( .A(n1381), .B(n1404), .CI(n1379), .CO(n1376), .S(n1377) );
  FA_X1 U1058 ( .A(n1383), .B(n1408), .CI(n1406), .CO(n1378), .S(n1379) );
  FA_X1 U1059 ( .A(n1410), .B(n1387), .CI(n1385), .CO(n1380), .S(n1381) );
  FA_X1 U1060 ( .A(n1389), .B(n1391), .CI(n1412), .CO(n1382), .S(n1383) );
  FA_X1 U1061 ( .A(n1416), .B(n1418), .CI(n1414), .CO(n1384), .S(n1385) );
  FA_X1 U1062 ( .A(n1399), .B(n1397), .CI(n1393), .CO(n1386), .S(n1387) );
  FA_X1 U1063 ( .A(n1401), .B(n1422), .CI(n1395), .CO(n1388), .S(n1389) );
  FA_X1 U1064 ( .A(n1420), .B(n1426), .CI(n1424), .CO(n1390), .S(n1391) );
  FA_X1 U1065 ( .A(n2438), .B(n2470), .CI(n2502), .CO(n1392), .S(n1393) );
  FA_X1 U1066 ( .A(n2406), .B(n2374), .CI(n2246), .CO(n1394), .S(n1395) );
  FA_X1 U1067 ( .A(n2118), .B(n2310), .CI(n2214), .CO(n1396), .S(n1397) );
  FA_X1 U1068 ( .A(n2150), .B(n2278), .CI(n2182), .CO(n1398), .S(n1399) );
  FA_X1 U1069 ( .A(n2089), .B(n1428), .CI(n2342), .CO(n1400), .S(n1401) );
  FA_X1 U1070 ( .A(n1432), .B(n1407), .CI(n1405), .CO(n1402), .S(n1403) );
  FA_X1 U1071 ( .A(n1409), .B(n1436), .CI(n1434), .CO(n1404), .S(n1405) );
  FA_X1 U1072 ( .A(n1438), .B(n1413), .CI(n1411), .CO(n1406), .S(n1407) );
  FA_X1 U1073 ( .A(n1415), .B(n1417), .CI(n1440), .CO(n1408), .S(n1409) );
  FA_X1 U1074 ( .A(n1419), .B(n1444), .CI(n1442), .CO(n1410), .S(n1411) );
  FA_X1 U1075 ( .A(n1425), .B(n1423), .CI(n1446), .CO(n1412), .S(n1413) );
  FA_X1 U1076 ( .A(n1427), .B(n1452), .CI(n1421), .CO(n1414), .S(n1415) );
  FA_X1 U1077 ( .A(n1448), .B(n1454), .CI(n1450), .CO(n1416), .S(n1417) );
  FA_X1 U1078 ( .A(n2247), .B(n2311), .CI(n1456), .CO(n1418), .S(n1419) );
  FA_X1 U1079 ( .A(n2183), .B(n2343), .CI(n2215), .CO(n1420), .S(n1421) );
  FA_X1 U1080 ( .A(n2151), .B(n2407), .CI(n2375), .CO(n1422), .S(n1423) );
  FA_X1 U1082 ( .A(n2503), .B(n1429), .CI(n2471), .CO(n1426), .S(n1427) );
  FA_X1 U1085 ( .A(n1437), .B(n1464), .CI(n1462), .CO(n1432), .S(n1433) );
  FA_X1 U1086 ( .A(n1466), .B(n1441), .CI(n1439), .CO(n1434), .S(n1435) );
  FA_X1 U1087 ( .A(n1443), .B(n1445), .CI(n1468), .CO(n1436), .S(n1437) );
  FA_X1 U1088 ( .A(n1472), .B(n1447), .CI(n1470), .CO(n1438), .S(n1439) );
  FA_X1 U1089 ( .A(n1453), .B(n1455), .CI(n1474), .CO(n1440), .S(n1441) );
  FA_X1 U1091 ( .A(n1482), .B(n1478), .CI(n1480), .CO(n1444), .S(n1445) );
  FA_X1 U1092 ( .A(n2536), .B(n1484), .CI(n1476), .CO(n1446), .S(n1447) );
  FA_X1 U1093 ( .A(n2280), .B(n2472), .CI(n2504), .CO(n1448), .S(n1449) );
  FA_X1 U1095 ( .A(n2152), .B(n2376), .CI(n2216), .CO(n1452), .S(n1453) );
  FA_X1 U1096 ( .A(n2120), .B(n2312), .CI(n2184), .CO(n1454), .S(n1455) );
  FA_X1 U1097 ( .A(n2090), .B(n1486), .CI(n2344), .CO(n1456), .S(n1457) );
  FA_X1 U1098 ( .A(n1490), .B(n1463), .CI(n1461), .CO(n1458), .S(n1459) );
  FA_X1 U1099 ( .A(n1465), .B(n1494), .CI(n1492), .CO(n1460), .S(n1461) );
  FA_X1 U1100 ( .A(n1496), .B(n1469), .CI(n1467), .CO(n1462), .S(n1463) );
  FA_X1 U1101 ( .A(n1471), .B(n1473), .CI(n1498), .CO(n1464), .S(n1465) );
  FA_X1 U1102 ( .A(n1500), .B(n1502), .CI(n1475), .CO(n1466), .S(n1467) );
  FA_X1 U1103 ( .A(n1506), .B(n1481), .CI(n1504), .CO(n1468), .S(n1469) );
  FA_X1 U1104 ( .A(n1483), .B(n1477), .CI(n1479), .CO(n1470), .S(n1471) );
  FA_X1 U1105 ( .A(n1514), .B(n1512), .CI(n1485), .CO(n1472), .S(n1473) );
  FA_X1 U1106 ( .A(n1508), .B(n1516), .CI(n1510), .CO(n1474), .S(n1475) );
  FA_X1 U1107 ( .A(n2249), .B(n2345), .CI(n2313), .CO(n1476), .S(n1477) );
  FA_X1 U1108 ( .A(n2185), .B(n2377), .CI(n2217), .CO(n1478), .S(n1479) );
  FA_X1 U1109 ( .A(n2441), .B(n2153), .CI(n2409), .CO(n1480), .S(n1481) );
  FA_X1 U1110 ( .A(n2473), .B(n2281), .CI(n2121), .CO(n1482), .S(n1483) );
  FA_X1 U1111 ( .A(n2537), .B(n1487), .CI(n2505), .CO(n1484), .S(n1485) );
  FA_X1 U1114 ( .A(n1495), .B(n1524), .CI(n1522), .CO(n1490), .S(n1491) );
  FA_X1 U1115 ( .A(n1499), .B(n1526), .CI(n1497), .CO(n1492), .S(n1493) );
  FA_X1 U1116 ( .A(n1501), .B(n1503), .CI(n1528), .CO(n1494), .S(n1495) );
  FA_X1 U1117 ( .A(n1532), .B(n1505), .CI(n1530), .CO(n1496), .S(n1497) );
  FA_X1 U1118 ( .A(n1534), .B(n1536), .CI(n1507), .CO(n1498), .S(n1499) );
  FA_X1 U1120 ( .A(n1517), .B(n1540), .CI(n1509), .CO(n1502), .S(n1503) );
  FA_X1 U1121 ( .A(n1544), .B(n1538), .CI(n1542), .CO(n1504), .S(n1505) );
  FA_X1 U1122 ( .A(n2570), .B(n2474), .CI(n1546), .CO(n1506), .S(n1507) );
  FA_X1 U1123 ( .A(n2506), .B(n2538), .CI(n2442), .CO(n1508), .S(n1509) );
  FA_X1 U1124 ( .A(n2346), .B(n2250), .CI(n2282), .CO(n1510), .S(n1511) );
  FA_X1 U1126 ( .A(n2154), .B(n2314), .CI(n2122), .CO(n1514), .S(n1515) );
  FA_X1 U1127 ( .A(n2091), .B(n1548), .CI(n2378), .CO(n1516), .S(n1517) );
  FA_X1 U1128 ( .A(n1552), .B(n1523), .CI(n1521), .CO(n1518), .S(n1519) );
  FA_X1 U1130 ( .A(n1529), .B(n1558), .CI(n1527), .CO(n1522), .S(n1523) );
  FA_X1 U1131 ( .A(n1531), .B(n1533), .CI(n1560), .CO(n1524), .S(n1525) );
  FA_X1 U1132 ( .A(n1562), .B(n1537), .CI(n1535), .CO(n1526), .S(n1527) );
  FA_X1 U1133 ( .A(n1566), .B(n1568), .CI(n1564), .CO(n1528), .S(n1529) );
  FA_X1 U1134 ( .A(n1543), .B(n1545), .CI(n1541), .CO(n1530), .S(n1531) );
  FA_X1 U1136 ( .A(n1576), .B(n1570), .CI(n1574), .CO(n1534), .S(n1535) );
  FA_X1 U1137 ( .A(n2411), .B(n2379), .CI(n1578), .CO(n1536), .S(n1537) );
  FA_X1 U1139 ( .A(n2475), .B(n2251), .CI(n2283), .CO(n1540), .S(n1541) );
  FA_X1 U1140 ( .A(n2187), .B(n2507), .CI(n2219), .CO(n1542), .S(n1543) );
  FA_X1 U1141 ( .A(n2155), .B(n2539), .CI(n2123), .CO(n1544), .S(n1545) );
  FA_X1 U1142 ( .A(n1580), .B(n2092), .CI(n2571), .CO(n1546), .S(n1547) );
  FA_X1 U1145 ( .A(n1557), .B(n1559), .CI(n1585), .CO(n1552), .S(n1553) );
  FA_X1 U1146 ( .A(n1561), .B(n1589), .CI(n1587), .CO(n1554), .S(n1555) );
  FA_X1 U1147 ( .A(n1591), .B(n1565), .CI(n1563), .CO(n1556), .S(n1557) );
  FA_X1 U1148 ( .A(n1593), .B(n1569), .CI(n1567), .CO(n1558), .S(n1559) );
  FA_X1 U1149 ( .A(n1597), .B(n1575), .CI(n1595), .CO(n1560), .S(n1561) );
  FA_X1 U1151 ( .A(n1599), .B(n1605), .CI(n1579), .CO(n1564), .S(n1565) );
  FA_X1 U1152 ( .A(n1607), .B(n1601), .CI(n1603), .CO(n1566), .S(n1567) );
  FA_X1 U1153 ( .A(n2604), .B(n2508), .CI(n1609), .CO(n1568), .S(n1569) );
  FA_X1 U1155 ( .A(n2284), .B(n2380), .CI(n2316), .CO(n1572), .S(n1573) );
  FA_X1 U1156 ( .A(n2252), .B(n2444), .CI(n2220), .CO(n1574), .S(n1575) );
  FA_X1 U1158 ( .A(n2412), .B(n1580), .CI(n2156), .CO(n1578), .S(n1579) );
  FA_X1 U1160 ( .A(n1613), .B(n1586), .CI(n1584), .CO(n1581), .S(n1582) );
  FA_X1 U1161 ( .A(n1588), .B(n1590), .CI(n1615), .CO(n1583), .S(n1584) );
  FA_X1 U1162 ( .A(n1619), .B(n1592), .CI(n1617), .CO(n1585), .S(n1586) );
  FA_X1 U1163 ( .A(n1621), .B(n1596), .CI(n1594), .CO(n1587), .S(n1588) );
  FA_X1 U1164 ( .A(n1623), .B(n1625), .CI(n1598), .CO(n1589), .S(n1590) );
  FA_X1 U1165 ( .A(n1600), .B(n1606), .CI(n1627), .CO(n1591), .S(n1592) );
  FA_X1 U1166 ( .A(n1608), .B(n1602), .CI(n1604), .CO(n1593), .S(n1594) );
  FA_X1 U1167 ( .A(n1633), .B(n1629), .CI(n1610), .CO(n1595), .S(n1596) );
  FA_X1 U1168 ( .A(n1637), .B(n1631), .CI(n1635), .CO(n1597), .S(n1598) );
  FA_X1 U1169 ( .A(n2445), .B(n2413), .CI(n1639), .CO(n1599), .S(n1600) );
  FA_X1 U1170 ( .A(n2317), .B(n2477), .CI(n2349), .CO(n1601), .S(n1602) );
  FA_X1 U1171 ( .A(n2253), .B(n2509), .CI(n2285), .CO(n1603), .S(n1604) );
  FA_X1 U1172 ( .A(n2541), .B(n2381), .CI(n2221), .CO(n1605), .S(n1606) );
  FA_X1 U1173 ( .A(n2125), .B(n2189), .CI(n2573), .CO(n1607), .S(n1608) );
  FA_X1 U1174 ( .A(n2157), .B(n2093), .CI(n2605), .CO(n1609), .S(n1610) );
  FA_X1 U1175 ( .A(n1643), .B(n1616), .CI(n1614), .CO(n1611), .S(n1612) );
  FA_X1 U1177 ( .A(n1649), .B(n1622), .CI(n1647), .CO(n1615), .S(n1616) );
  FA_X1 U1178 ( .A(n1651), .B(n1626), .CI(n1624), .CO(n1617), .S(n1618) );
  FA_X1 U1179 ( .A(n1628), .B(n1655), .CI(n1653), .CO(n1619), .S(n1620) );
  FA_X1 U1180 ( .A(n1632), .B(n1634), .CI(n1657), .CO(n1621), .S(n1622) );
  FA_X1 U1181 ( .A(n1638), .B(n1630), .CI(n1636), .CO(n1623), .S(n1624) );
  FA_X1 U1182 ( .A(n1663), .B(n1659), .CI(n1661), .CO(n1625), .S(n1626) );
  FA_X1 U1183 ( .A(n1667), .B(n1640), .CI(n1665), .CO(n1627), .S(n1628) );
  FA_X1 U1184 ( .A(n2414), .B(n2286), .CI(n2350), .CO(n1629), .S(n1630) );
  FA_X1 U1185 ( .A(n2190), .B(n2446), .CI(n2222), .CO(n1631), .S(n1632) );
  FA_X1 U1186 ( .A(n2158), .B(n2254), .CI(n2478), .CO(n1633), .S(n1634) );
  FA_X1 U1187 ( .A(n2542), .B(n2318), .CI(n2510), .CO(n1635), .S(n1636) );
  FA_X1 U1188 ( .A(n2574), .B(n2382), .CI(n2606), .CO(n1637), .S(n1638) );
  HA_X1 U1189 ( .A(n2061), .B(n2126), .CO(n1639), .S(n1640) );
  FA_X1 U1190 ( .A(n1671), .B(n1646), .CI(n1644), .CO(n1641), .S(n1642) );
  FA_X1 U1191 ( .A(n1648), .B(n1650), .CI(n1673), .CO(n1643), .S(n1644) );
  FA_X1 U1192 ( .A(n1677), .B(n1652), .CI(n1675), .CO(n1645), .S(n1646) );
  FA_X1 U1193 ( .A(n1656), .B(n1679), .CI(n1654), .CO(n1647), .S(n1648) );
  FA_X1 U1194 ( .A(n1681), .B(n1683), .CI(n1658), .CO(n1649), .S(n1650) );
  FA_X1 U1195 ( .A(n1664), .B(n1662), .CI(n1685), .CO(n1651), .S(n1652) );
  FA_X1 U1196 ( .A(n1668), .B(n1660), .CI(n1666), .CO(n1653), .S(n1654) );
  FA_X1 U1197 ( .A(n1691), .B(n1687), .CI(n1689), .CO(n1655), .S(n1656) );
  FA_X1 U1198 ( .A(n1695), .B(n2447), .CI(n1693), .CO(n1657), .S(n1658) );
  FA_X1 U1199 ( .A(n2479), .B(n2383), .CI(n2415), .CO(n1659), .S(n1660) );
  FA_X1 U1200 ( .A(n2319), .B(n2287), .CI(n2351), .CO(n1661), .S(n1662) );
  FA_X1 U1201 ( .A(n2223), .B(n2511), .CI(n2255), .CO(n1663), .S(n1664) );
  FA_X1 U1202 ( .A(n2191), .B(n2575), .CI(n2543), .CO(n1665), .S(n1666) );
  FA_X1 U1203 ( .A(n2159), .B(n2607), .CI(n2127), .CO(n1667), .S(n1668) );
  FA_X1 U1205 ( .A(n1676), .B(n1678), .CI(n1701), .CO(n1671), .S(n1672) );
  FA_X1 U1206 ( .A(n1705), .B(n1680), .CI(n1703), .CO(n1673), .S(n1674) );
  FA_X1 U1207 ( .A(n1684), .B(n1707), .CI(n1682), .CO(n1675), .S(n1676) );
  FA_X1 U1208 ( .A(n1686), .B(n1711), .CI(n1709), .CO(n1677), .S(n1678) );
  FA_X1 U1209 ( .A(n1690), .B(n1692), .CI(n1694), .CO(n1679), .S(n1680) );
  FA_X1 U1210 ( .A(n1713), .B(n1717), .CI(n1688), .CO(n1681), .S(n1682) );
  FA_X1 U1211 ( .A(n1721), .B(n1715), .CI(n1719), .CO(n1683), .S(n1684) );
  FA_X1 U1212 ( .A(n2480), .B(n2448), .CI(n1696), .CO(n1685), .S(n1686) );
  FA_X1 U1213 ( .A(n2288), .B(n2512), .CI(n2320), .CO(n1687), .S(n1688) );
  FA_X1 U1214 ( .A(n2544), .B(n2416), .CI(n2256), .CO(n1689), .S(n1690) );
  FA_X1 U1215 ( .A(n2576), .B(n2352), .CI(n2224), .CO(n1691), .S(n1692) );
  FA_X1 U1216 ( .A(n2608), .B(n2192), .CI(n2384), .CO(n1693), .S(n1694) );
  HA_X1 U1217 ( .A(n2160), .B(n2062), .CO(n1695), .S(n1696) );
  FA_X1 U1218 ( .A(n1725), .B(n1702), .CI(n1700), .CO(n1697), .S(n1698) );
  FA_X1 U1219 ( .A(n1704), .B(n1729), .CI(n1727), .CO(n1699), .S(n1700) );
  FA_X1 U1220 ( .A(n1731), .B(n1708), .CI(n1706), .CO(n1701), .S(n1702) );
  FA_X1 U1221 ( .A(n1733), .B(n1712), .CI(n1710), .CO(n1703), .S(n1704) );
  FA_X1 U1222 ( .A(n1737), .B(n1718), .CI(n1735), .CO(n1705), .S(n1706) );
  FA_X1 U1223 ( .A(n1722), .B(n1716), .CI(n1720), .CO(n1707), .S(n1708) );
  FA_X1 U1224 ( .A(n1741), .B(n1739), .CI(n1714), .CO(n1709), .S(n1710) );
  FA_X1 U1225 ( .A(n1745), .B(n1747), .CI(n1743), .CO(n1711), .S(n1712) );
  FA_X1 U1226 ( .A(n2417), .B(n2385), .CI(n2449), .CO(n1713), .S(n1714) );
  FA_X1 U1227 ( .A(n2321), .B(n2481), .CI(n2353), .CO(n1715), .S(n1716) );
  FA_X1 U1228 ( .A(n2257), .B(n2513), .CI(n2289), .CO(n1717), .S(n1718) );
  FA_X1 U1229 ( .A(n2225), .B(n2577), .CI(n2545), .CO(n1719), .S(n1720) );
  FA_X1 U1230 ( .A(n2193), .B(n2609), .CI(n2161), .CO(n1721), .S(n1722) );
  FA_X1 U1232 ( .A(n1730), .B(n1732), .CI(n1753), .CO(n1725), .S(n1726) );
  FA_X1 U1233 ( .A(n1734), .B(n1757), .CI(n1755), .CO(n1727), .S(n1728) );
  FA_X1 U1234 ( .A(n1759), .B(n1738), .CI(n1736), .CO(n1729), .S(n1730) );
  FA_X1 U1235 ( .A(n1744), .B(n1746), .CI(n1761), .CO(n1731), .S(n1732) );
  FA_X1 U1236 ( .A(n1740), .B(n1763), .CI(n1742), .CO(n1733), .S(n1734) );
  FA_X1 U1237 ( .A(n1767), .B(n1765), .CI(n1769), .CO(n1735), .S(n1736) );
  FA_X1 U1238 ( .A(n1748), .B(n2514), .CI(n1771), .CO(n1737), .S(n1738) );
  FA_X1 U1240 ( .A(n2578), .B(n2354), .CI(n2322), .CO(n1741), .S(n1742) );
  FA_X1 U1241 ( .A(n2258), .B(n2386), .CI(n2290), .CO(n1743), .S(n1744) );
  FA_X1 U1242 ( .A(n2610), .B(n2418), .CI(n2226), .CO(n1745), .S(n1746) );
  HA_X1 U1243 ( .A(n2194), .B(n2063), .CO(n1747), .S(n1748) );
  FA_X1 U1245 ( .A(n1777), .B(n1779), .CI(n1756), .CO(n1751), .S(n1752) );
  FA_X1 U1246 ( .A(n1760), .B(n1762), .CI(n1758), .CO(n1753), .S(n1754) );
  FA_X1 U1247 ( .A(n1783), .B(n1785), .CI(n1781), .CO(n1755), .S(n1756) );
  FA_X1 U1248 ( .A(n1770), .B(n1772), .CI(n1764), .CO(n1757), .S(n1758) );
  FA_X1 U1249 ( .A(n1766), .B(n1793), .CI(n1768), .CO(n1759), .S(n1760) );
  FA_X1 U1250 ( .A(n1787), .B(n1789), .CI(n1791), .CO(n1761), .S(n1762) );
  FA_X1 U1251 ( .A(n2451), .B(n2483), .CI(n1795), .CO(n1763), .S(n1764) );
  FA_X1 U1252 ( .A(n2387), .B(n2515), .CI(n2419), .CO(n1765), .S(n1766) );
  FA_X1 U1253 ( .A(n2355), .B(n2547), .CI(n2323), .CO(n1767), .S(n1768) );
  FA_X1 U1254 ( .A(n2259), .B(n2579), .CI(n2291), .CO(n1769), .S(n1770) );
  FA_X1 U1255 ( .A(n2195), .B(n2611), .CI(n2227), .CO(n1771), .S(n1772) );
  FA_X1 U1256 ( .A(n1799), .B(n1778), .CI(n1776), .CO(n1773), .S(n1774) );
  FA_X1 U1257 ( .A(n1803), .B(n1780), .CI(n1801), .CO(n1775), .S(n1776) );
  FA_X1 U1258 ( .A(n1784), .B(n1805), .CI(n1782), .CO(n1777), .S(n1778) );
  FA_X1 U1259 ( .A(n1807), .B(n1809), .CI(n1786), .CO(n1779), .S(n1780) );
  FA_X1 U1260 ( .A(n1794), .B(n1790), .CI(n1792), .CO(n1781), .S(n1782) );
  FA_X1 U1261 ( .A(n1811), .B(n1813), .CI(n1788), .CO(n1783), .S(n1784) );
  FA_X1 U1262 ( .A(n1817), .B(n1796), .CI(n1815), .CO(n1785), .S(n1786) );
  FA_X1 U1263 ( .A(n2356), .B(n2484), .CI(n2452), .CO(n1787), .S(n1788) );
  FA_X1 U1264 ( .A(n2292), .B(n2516), .CI(n2324), .CO(n1789), .S(n1790) );
  FA_X1 U1265 ( .A(n2580), .B(n2388), .CI(n2548), .CO(n1791), .S(n1792) );
  FA_X1 U1266 ( .A(n2612), .B(n2260), .CI(n2420), .CO(n1793), .S(n1794) );
  HA_X1 U1267 ( .A(n2228), .B(n2064), .CO(n1795), .S(n1796) );
  FA_X1 U1268 ( .A(n1821), .B(n1802), .CI(n1800), .CO(n1797), .S(n1798) );
  FA_X1 U1269 ( .A(n1804), .B(n1825), .CI(n1823), .CO(n1799), .S(n1800) );
  FA_X1 U1270 ( .A(n1808), .B(n1827), .CI(n1806), .CO(n1801), .S(n1802) );
  FA_X1 U1271 ( .A(n1829), .B(n1831), .CI(n1810), .CO(n1803), .S(n1804) );
  FA_X1 U1272 ( .A(n1818), .B(n1814), .CI(n1816), .CO(n1805), .S(n1806) );
  FA_X1 U1273 ( .A(n1833), .B(n1835), .CI(n1812), .CO(n1807), .S(n1808) );
  FA_X1 U1274 ( .A(n1839), .B(n2453), .CI(n1837), .CO(n1809), .S(n1810) );
  FA_X1 U1275 ( .A(n2485), .B(n2389), .CI(n2421), .CO(n1811), .S(n1812) );
  FA_X1 U1276 ( .A(n2357), .B(n2549), .CI(n2517), .CO(n1813), .S(n1814) );
  FA_X1 U1277 ( .A(n2293), .B(n2581), .CI(n2325), .CO(n1815), .S(n1816) );
  FA_X1 U1278 ( .A(n2261), .B(n2613), .CI(n2229), .CO(n1817), .S(n1818) );
  FA_X1 U1279 ( .A(n1843), .B(n1824), .CI(n1822), .CO(n1819), .S(n1820) );
  FA_X1 U1280 ( .A(n1845), .B(n1828), .CI(n1826), .CO(n1821), .S(n1822) );
  FA_X1 U1281 ( .A(n1830), .B(n1849), .CI(n1847), .CO(n1823), .S(n1824) );
  FA_X1 U1282 ( .A(n1851), .B(n1838), .CI(n1832), .CO(n1825), .S(n1826) );
  FA_X1 U1283 ( .A(n1834), .B(n1857), .CI(n1836), .CO(n1827), .S(n1828) );
  FA_X1 U1284 ( .A(n1853), .B(n1859), .CI(n1855), .CO(n1829), .S(n1830) );
  FA_X1 U1285 ( .A(n2486), .B(n2518), .CI(n1840), .CO(n1831), .S(n1832) );
  FA_X1 U1286 ( .A(n2358), .B(n2550), .CI(n2390), .CO(n1833), .S(n1834) );
  FA_X1 U1287 ( .A(n2582), .B(n2422), .CI(n2326), .CO(n1835), .S(n1836) );
  FA_X1 U1288 ( .A(n2614), .B(n2454), .CI(n2294), .CO(n1837), .S(n1838) );
  HA_X1 U1289 ( .A(n2262), .B(n2065), .CO(n1839), .S(n1840) );
  FA_X1 U1290 ( .A(n1863), .B(n1846), .CI(n1844), .CO(n1841), .S(n1842) );
  FA_X1 U1291 ( .A(n1848), .B(n1850), .CI(n1865), .CO(n1843), .S(n1844) );
  FA_X1 U1293 ( .A(n1860), .B(n1858), .CI(n1871), .CO(n1847), .S(n1848) );
  FA_X1 U1294 ( .A(n1854), .B(n1873), .CI(n1856), .CO(n1849), .S(n1850) );
  FA_X1 U1297 ( .A(n2391), .B(n2551), .CI(n2423), .CO(n1855), .S(n1856) );
  FA_X1 U1298 ( .A(n2327), .B(n2583), .CI(n2359), .CO(n1857), .S(n1858) );
  FA_X1 U1299 ( .A(n2295), .B(n2615), .CI(n2263), .CO(n1859), .S(n1860) );
  FA_X1 U1300 ( .A(n1883), .B(n1866), .CI(n1864), .CO(n1861), .S(n1862) );
  FA_X1 U1301 ( .A(n1868), .B(n1870), .CI(n1885), .CO(n1863), .S(n1864) );
  FA_X1 U1302 ( .A(n1872), .B(n1889), .CI(n1887), .CO(n1865), .S(n1866) );
  FA_X1 U1303 ( .A(n1878), .B(n1874), .CI(n1876), .CO(n1867), .S(n1868) );
  FA_X1 U1304 ( .A(n1893), .B(n1895), .CI(n1891), .CO(n1869), .S(n1870) );
  FA_X1 U1305 ( .A(n1880), .B(n2488), .CI(n1897), .CO(n1871), .S(n1872) );
  FA_X1 U1306 ( .A(n2360), .B(n2520), .CI(n2392), .CO(n1873), .S(n1874) );
  FA_X1 U1307 ( .A(n2328), .B(n2424), .CI(n2552), .CO(n1875), .S(n1876) );
  FA_X1 U1308 ( .A(n2616), .B(n2456), .CI(n2584), .CO(n1877), .S(n1878) );
  HA_X1 U1309 ( .A(n2296), .B(n2066), .CO(n1879), .S(n1880) );
  FA_X1 U1310 ( .A(n1901), .B(n1886), .CI(n1884), .CO(n1881), .S(n1882) );
  FA_X1 U1311 ( .A(n1888), .B(n1890), .CI(n1903), .CO(n1883), .S(n1884) );
  FA_X1 U1312 ( .A(n1907), .B(n1892), .CI(n1905), .CO(n1885), .S(n1886) );
  FA_X1 U1313 ( .A(n1898), .B(n1894), .CI(n1896), .CO(n1887), .S(n1888) );
  FA_X1 U1314 ( .A(n1909), .B(n1913), .CI(n1911), .CO(n1889), .S(n1890) );
  FA_X1 U1315 ( .A(n2489), .B(n2521), .CI(n1915), .CO(n1891), .S(n1892) );
  FA_X1 U1316 ( .A(n2425), .B(n2553), .CI(n2457), .CO(n1893), .S(n1894) );
  FA_X1 U1317 ( .A(n2361), .B(n2585), .CI(n2393), .CO(n1895), .S(n1896) );
  FA_X1 U1318 ( .A(n2329), .B(n2617), .CI(n2297), .CO(n1897), .S(n1898) );
  FA_X1 U1319 ( .A(n1919), .B(n1904), .CI(n1902), .CO(n1899), .S(n1900) );
  FA_X1 U1320 ( .A(n1906), .B(n1923), .CI(n1921), .CO(n1901), .S(n1902) );
  FA_X1 U1321 ( .A(n1925), .B(n1914), .CI(n1908), .CO(n1903), .S(n1904) );
  FA_X1 U1323 ( .A(n1931), .B(n1916), .CI(n1929), .CO(n1907), .S(n1908) );
  FA_X1 U1325 ( .A(n2618), .B(n2522), .CI(n2426), .CO(n1911), .S(n1912) );
  FA_X1 U1326 ( .A(n2362), .B(n2490), .CI(n2394), .CO(n1913), .S(n1914) );
  HA_X1 U1327 ( .A(n2330), .B(n2067), .CO(n1915), .S(n1916) );
  FA_X1 U1328 ( .A(n1935), .B(n1922), .CI(n1920), .CO(n1917), .S(n1918) );
  FA_X1 U1329 ( .A(n1924), .B(n1926), .CI(n1937), .CO(n1919), .S(n1920) );
  FA_X1 U1330 ( .A(n1941), .B(n1932), .CI(n1939), .CO(n1921), .S(n1922) );
  FA_X1 U1331 ( .A(n1928), .B(n1943), .CI(n1930), .CO(n1923), .S(n1924) );
  FA_X1 U1332 ( .A(n1947), .B(n2523), .CI(n1945), .CO(n1925), .S(n1926) );
  FA_X1 U1333 ( .A(n2459), .B(n2555), .CI(n2491), .CO(n1927), .S(n1928) );
  FA_X1 U1334 ( .A(n2395), .B(n2587), .CI(n2427), .CO(n1929), .S(n1930) );
  FA_X1 U1335 ( .A(n2363), .B(n2619), .CI(n2331), .CO(n1931), .S(n1932) );
  FA_X1 U1336 ( .A(n1938), .B(n1951), .CI(n1936), .CO(n1933), .S(n1934) );
  FA_X1 U1337 ( .A(n1953), .B(n1942), .CI(n1940), .CO(n1935), .S(n1936) );
  FA_X1 U1338 ( .A(n1946), .B(n1944), .CI(n1955), .CO(n1937), .S(n1938) );
  FA_X1 U1339 ( .A(n1957), .B(n1961), .CI(n1959), .CO(n1939), .S(n1940) );
  FA_X1 U1340 ( .A(n2556), .B(n2588), .CI(n1948), .CO(n1941), .S(n1942) );
  FA_X1 U1341 ( .A(n2428), .B(n2524), .CI(n2460), .CO(n1943), .S(n1944) );
  FA_X1 U1342 ( .A(n2396), .B(n2492), .CI(n2620), .CO(n1945), .S(n1946) );
  HA_X1 U1343 ( .A(n2364), .B(n2068), .CO(n1947), .S(n1948) );
  FA_X1 U1344 ( .A(n1965), .B(n1954), .CI(n1952), .CO(n1949), .S(n1950) );
  FA_X1 U1345 ( .A(n1967), .B(n1969), .CI(n1956), .CO(n1951), .S(n1952) );
  FA_X1 U1346 ( .A(n1960), .B(n1962), .CI(n1958), .CO(n1953), .S(n1954) );
  FA_X1 U1347 ( .A(n1973), .B(n1975), .CI(n1971), .CO(n1955), .S(n1956) );
  FA_X1 U1348 ( .A(n2493), .B(n2557), .CI(n2525), .CO(n1957), .S(n1958) );
  FA_X1 U1349 ( .A(n2429), .B(n2589), .CI(n2461), .CO(n1959), .S(n1960) );
  FA_X1 U1350 ( .A(n2397), .B(n2621), .CI(n2365), .CO(n1961), .S(n1962) );
  FA_X1 U1351 ( .A(n1979), .B(n1968), .CI(n1966), .CO(n1963), .S(n1964) );
  FA_X1 U1352 ( .A(n1981), .B(n1974), .CI(n1970), .CO(n1965), .S(n1966) );
  FA_X1 U1353 ( .A(n1983), .B(n1985), .CI(n1972), .CO(n1967), .S(n1968) );
  FA_X1 U1354 ( .A(n1976), .B(n2494), .CI(n1987), .CO(n1969), .S(n1970) );
  FA_X1 U1355 ( .A(n2558), .B(n2430), .CI(n2462), .CO(n1971), .S(n1972) );
  FA_X1 U1356 ( .A(n2622), .B(n2526), .CI(n2590), .CO(n1973), .S(n1974) );
  HA_X1 U1357 ( .A(n2398), .B(n2069), .CO(n1975), .S(n1976) );
  FA_X1 U1358 ( .A(n1991), .B(n1982), .CI(n1980), .CO(n1977), .S(n1978) );
  FA_X1 U1359 ( .A(n1984), .B(n1988), .CI(n1993), .CO(n1979), .S(n1980) );
  FA_X1 U1360 ( .A(n1995), .B(n1997), .CI(n1986), .CO(n1981), .S(n1982) );
  FA_X1 U1361 ( .A(n2527), .B(n2559), .CI(n1999), .CO(n1983), .S(n1984) );
  FA_X1 U1362 ( .A(n2463), .B(n2591), .CI(n2495), .CO(n1985), .S(n1986) );
  FA_X1 U1363 ( .A(n2431), .B(n2623), .CI(n2399), .CO(n1987), .S(n1988) );
  FA_X1 U1364 ( .A(n2003), .B(n1994), .CI(n1992), .CO(n1989), .S(n1990) );
  FA_X1 U1365 ( .A(n1998), .B(n1996), .CI(n2005), .CO(n1991), .S(n1992) );
  FA_X1 U1366 ( .A(n2009), .B(n2000), .CI(n2007), .CO(n1993), .S(n1994) );
  FA_X1 U1367 ( .A(n2464), .B(n2560), .CI(n2496), .CO(n1995), .S(n1996) );
  FA_X1 U1368 ( .A(n2624), .B(n2528), .CI(n2592), .CO(n1997), .S(n1998) );
  HA_X1 U1369 ( .A(n2432), .B(n2070), .CO(n1999), .S(n2000) );
  FA_X1 U1370 ( .A(n2006), .B(n2013), .CI(n2004), .CO(n2001), .S(n2002) );
  FA_X1 U1371 ( .A(n2010), .B(n2008), .CI(n2015), .CO(n2003), .S(n2004) );
  FA_X1 U1372 ( .A(n2019), .B(n2561), .CI(n2017), .CO(n2005), .S(n2006) );
  FA_X1 U1373 ( .A(n2497), .B(n2593), .CI(n2529), .CO(n2007), .S(n2008) );
  FA_X1 U1374 ( .A(n2465), .B(n2625), .CI(n2433), .CO(n2009), .S(n2010) );
  FA_X1 U1375 ( .A(n2023), .B(n2016), .CI(n2014), .CO(n2011), .S(n2012) );
  FA_X1 U1376 ( .A(n2025), .B(n2027), .CI(n2018), .CO(n2013), .S(n2014) );
  FA_X1 U1377 ( .A(n2498), .B(n2530), .CI(n2020), .CO(n2015), .S(n2016) );
  FA_X1 U1378 ( .A(n2626), .B(n2562), .CI(n2594), .CO(n2017), .S(n2018) );
  HA_X1 U1379 ( .A(n2466), .B(n2071), .CO(n2019), .S(n2020) );
  FA_X1 U1380 ( .A(n2031), .B(n2028), .CI(n2024), .CO(n2021), .S(n2022) );
  FA_X1 U1381 ( .A(n2033), .B(n2035), .CI(n2026), .CO(n2023), .S(n2024) );
  FA_X1 U1382 ( .A(n2531), .B(n2595), .CI(n2563), .CO(n2025), .S(n2026) );
  FA_X1 U1383 ( .A(n2499), .B(n2627), .CI(n2467), .CO(n2027), .S(n2028) );
  FA_X1 U1384 ( .A(n2034), .B(n2039), .CI(n2032), .CO(n2029), .S(n2030) );
  FA_X1 U1385 ( .A(n2036), .B(n2628), .CI(n2041), .CO(n2031), .S(n2032) );
  FA_X1 U1386 ( .A(n2532), .B(n2564), .CI(n2596), .CO(n2033), .S(n2034) );
  HA_X1 U1387 ( .A(n2500), .B(n2072), .CO(n2035), .S(n2036) );
  FA_X1 U1388 ( .A(n2042), .B(n2045), .CI(n2040), .CO(n2037), .S(n2038) );
  FA_X1 U1389 ( .A(n2565), .B(n2597), .CI(n2047), .CO(n2039), .S(n2040) );
  FA_X1 U1390 ( .A(n2533), .B(n2629), .CI(n2501), .CO(n2041), .S(n2042) );
  FA_X1 U1391 ( .A(n2051), .B(n2048), .CI(n2046), .CO(n2043), .S(n2044) );
  FA_X1 U1392 ( .A(n2566), .B(n2630), .CI(n2598), .CO(n2045), .S(n2046) );
  HA_X1 U1393 ( .A(n2534), .B(n2073), .CO(n2047), .S(n2048) );
  FA_X1 U1394 ( .A(n2055), .B(n2599), .CI(n2052), .CO(n2049), .S(n2050) );
  FA_X1 U1395 ( .A(n2567), .B(n2631), .CI(n2535), .CO(n2051), .S(n2052) );
  FA_X1 U1396 ( .A(n2600), .B(n2632), .CI(n2056), .CO(n2053), .S(n2054) );
  HA_X1 U1397 ( .A(n2568), .B(n2074), .CO(n2055), .S(n2056) );
  FA_X1 U1398 ( .A(n2601), .B(n2633), .CI(n2569), .CO(n2057), .S(n2058) );
  HA_X1 U1399 ( .A(n2634), .B(n2602), .CO(n2059), .S(n2060) );
  NOR2_X4 U1400 ( .A1(n2637), .A2(n3462), .ZN(n2077) );
  NOR2_X4 U1401 ( .A1(n2638), .A2(n3462), .ZN(n1044) );
  NOR2_X4 U1402 ( .A1(n2639), .A2(n3462), .ZN(n2078) );
  NOR2_X4 U1403 ( .A1(n2640), .A2(n3462), .ZN(n1054) );
  NOR2_X4 U1404 ( .A1(n2641), .A2(n3462), .ZN(n2079) );
  NOR2_X4 U1405 ( .A1(n2642), .A2(n3462), .ZN(n1068) );
  NOR2_X4 U1406 ( .A1(n2643), .A2(n3462), .ZN(n2080) );
  NOR2_X4 U1407 ( .A1(n2644), .A2(n3462), .ZN(n1086) );
  NOR2_X4 U1408 ( .A1(n2645), .A2(n3462), .ZN(n2081) );
  NOR2_X4 U1409 ( .A1(n2646), .A2(n3462), .ZN(n1108) );
  NOR2_X4 U1410 ( .A1(n2647), .A2(n3462), .ZN(n2082) );
  NOR2_X4 U1411 ( .A1(n2648), .A2(n3462), .ZN(n1134) );
  NOR2_X4 U1412 ( .A1(n2649), .A2(n3462), .ZN(n2083) );
  NOR2_X4 U1413 ( .A1(n2650), .A2(n3462), .ZN(n1164) );
  NOR2_X4 U1414 ( .A1(n2651), .A2(n3462), .ZN(n2084) );
  NOR2_X4 U1415 ( .A1(n2652), .A2(n3462), .ZN(n1198) );
  NOR2_X4 U1416 ( .A1(n2653), .A2(n3462), .ZN(n2085) );
  NOR2_X4 U1417 ( .A1(n2654), .A2(n3462), .ZN(n1236) );
  NOR2_X4 U1418 ( .A1(n2655), .A2(n3462), .ZN(n2086) );
  NOR2_X4 U1419 ( .A1(n2656), .A2(n3462), .ZN(n1278) );
  NOR2_X4 U1420 ( .A1(n2657), .A2(n3462), .ZN(n2087) );
  NOR2_X4 U1421 ( .A1(n2658), .A2(n3462), .ZN(n1324) );
  NOR2_X4 U1422 ( .A1(n2659), .A2(n3462), .ZN(n2088) );
  NOR2_X4 U1423 ( .A1(n2660), .A2(n3462), .ZN(n1374) );
  NOR2_X4 U1424 ( .A1(n2661), .A2(n3462), .ZN(n2089) );
  NOR2_X4 U1426 ( .A1(n2663), .A2(n3462), .ZN(n2090) );
  NOR2_X4 U1428 ( .A1(n2665), .A2(n3462), .ZN(n2091) );
  NOR2_X4 U1429 ( .A1(n2666), .A2(n3462), .ZN(n2092) );
  NOR2_X4 U1430 ( .A1(n2667), .A2(n3462), .ZN(n1548) );
  OAI22_X2 U1463 ( .A1(n3663), .A2(n2668), .B1(n3654), .B2(n3462), .ZN(n2095)
         );
  OAI22_X2 U1464 ( .A1(n3663), .A2(n2669), .B1(n2668), .B2(n3655), .ZN(n2096)
         );
  OAI22_X2 U1465 ( .A1(n3663), .A2(n2670), .B1(n2669), .B2(n3654), .ZN(n2097)
         );
  OAI22_X2 U1466 ( .A1(n3663), .A2(n2671), .B1(n2670), .B2(n3654), .ZN(n2098)
         );
  OAI22_X2 U1467 ( .A1(n3663), .A2(n2672), .B1(n2671), .B2(n3655), .ZN(n2099)
         );
  OAI22_X2 U1469 ( .A1(n3663), .A2(n2674), .B1(n2673), .B2(n3655), .ZN(n2101)
         );
  OAI22_X2 U1594 ( .A1(n3729), .A2(n2735), .B1(n2734), .B2(n408), .ZN(n2164)
         );
  OAI22_X2 U1595 ( .A1(n3729), .A2(n2736), .B1(n2735), .B2(n408), .ZN(n2165)
         );
  OAI22_X2 U1596 ( .A1(n3729), .A2(n2737), .B1(n2736), .B2(n408), .ZN(n2166)
         );
  OAI22_X2 U1597 ( .A1(n3729), .A2(n2738), .B1(n2737), .B2(n408), .ZN(n2167)
         );
  OAI22_X2 U1599 ( .A1(n3729), .A2(n2740), .B1(n2739), .B2(n408), .ZN(n2169)
         );
  OAI22_X2 U1601 ( .A1(n3729), .A2(n2742), .B1(n2741), .B2(n408), .ZN(n2171)
         );
  OAI22_X2 U1602 ( .A1(n3729), .A2(n2743), .B1(n2742), .B2(n408), .ZN(n2172)
         );
  OAI22_X2 U1603 ( .A1(n3729), .A2(n2744), .B1(n2743), .B2(n408), .ZN(n2173)
         );
  OAI22_X2 U1658 ( .A1(n3471), .A2(n2767), .B1(n3631), .B2(n3730), .ZN(n2197)
         );
  OAI22_X2 U1659 ( .A1(n3471), .A2(n2768), .B1(n2767), .B2(n3630), .ZN(n2198)
         );
  OAI22_X2 U1660 ( .A1(n3471), .A2(n2769), .B1(n2768), .B2(n3631), .ZN(n2199)
         );
  OAI22_X2 U1661 ( .A1(n3471), .A2(n2770), .B1(n2769), .B2(n3631), .ZN(n2200)
         );
  OAI22_X2 U1662 ( .A1(n3471), .A2(n2771), .B1(n2770), .B2(n3631), .ZN(n2201)
         );
  OAI22_X2 U1663 ( .A1(n3471), .A2(n2772), .B1(n2771), .B2(n3630), .ZN(n2202)
         );
  OAI22_X2 U1664 ( .A1(n3471), .A2(n2773), .B1(n2772), .B2(n3630), .ZN(n2203)
         );
  OAI22_X2 U1665 ( .A1(n3471), .A2(n2774), .B1(n2773), .B2(n3631), .ZN(n2204)
         );
  OAI22_X2 U1666 ( .A1(n3471), .A2(n2775), .B1(n2774), .B2(n3630), .ZN(n2205)
         );
  OAI22_X2 U1668 ( .A1(n3471), .A2(n2777), .B1(n2776), .B2(n3630), .ZN(n2207)
         );
  OAI22_X2 U1669 ( .A1(n3471), .A2(n2778), .B1(n2777), .B2(n3631), .ZN(n2208)
         );
  OAI22_X2 U1670 ( .A1(n455), .A2(n2779), .B1(n2778), .B2(n3631), .ZN(n2209)
         );
  OAI22_X2 U1671 ( .A1(n455), .A2(n2780), .B1(n2779), .B2(n3630), .ZN(n2210)
         );
  OAI22_X2 U1672 ( .A1(n3471), .A2(n2781), .B1(n2780), .B2(n3631), .ZN(n2211)
         );
  OAI22_X2 U1673 ( .A1(n3471), .A2(n2782), .B1(n2781), .B2(n3631), .ZN(n2212)
         );
  OAI22_X2 U1674 ( .A1(n3471), .A2(n2783), .B1(n2782), .B2(n3631), .ZN(n2213)
         );
  OAI22_X2 U1676 ( .A1(n455), .A2(n2785), .B1(n2784), .B2(n3631), .ZN(n2215)
         );
  OAI22_X2 U1677 ( .A1(n3471), .A2(n2786), .B1(n2785), .B2(n3630), .ZN(n2216)
         );
  OAI22_X2 U1678 ( .A1(n455), .A2(n2787), .B1(n2786), .B2(n3631), .ZN(n2217)
         );
  OAI22_X2 U1681 ( .A1(n3471), .A2(n2790), .B1(n2789), .B2(n3630), .ZN(n2220)
         );
  OAI22_X2 U1682 ( .A1(n3471), .A2(n2791), .B1(n2790), .B2(n3630), .ZN(n2221)
         );
  OAI22_X2 U1683 ( .A1(n3471), .A2(n2792), .B1(n2791), .B2(n3630), .ZN(n2222)
         );
  OAI22_X2 U1684 ( .A1(n3471), .A2(n2793), .B1(n2792), .B2(n3630), .ZN(n2223)
         );
  OAI22_X2 U1685 ( .A1(n3471), .A2(n2794), .B1(n2793), .B2(n3631), .ZN(n2224)
         );
  OAI22_X2 U1686 ( .A1(n455), .A2(n2795), .B1(n2794), .B2(n3631), .ZN(n2225)
         );
  OAI22_X2 U1689 ( .A1(n455), .A2(n2798), .B1(n2797), .B2(n3631), .ZN(n2228)
         );
  OAI22_X2 U1728 ( .A1(n452), .A2(n2805), .B1(n2804), .B2(n402), .ZN(n2236) );
  OAI22_X2 U1735 ( .A1(n452), .A2(n2812), .B1(n2811), .B2(n402), .ZN(n2243) );
  OAI22_X2 U1742 ( .A1(n452), .A2(n2819), .B1(n2818), .B2(n402), .ZN(n2250) );
  OAI22_X2 U1753 ( .A1(n452), .A2(n2830), .B1(n2829), .B2(n402), .ZN(n2261) );
  OAI22_X2 U1787 ( .A1(n3475), .A2(n3282), .B1(n2865), .B2(n3672), .ZN(n2066)
         );
  OAI22_X2 U1788 ( .A1(n3474), .A2(n2833), .B1(n3672), .B2(n3282), .ZN(n2265)
         );
  OAI22_X2 U1789 ( .A1(n3474), .A2(n2834), .B1(n2833), .B2(n3673), .ZN(n2266)
         );
  OAI22_X2 U1790 ( .A1(n3475), .A2(n2835), .B1(n2834), .B2(n3673), .ZN(n2267)
         );
  OAI22_X2 U1791 ( .A1(n3474), .A2(n2836), .B1(n2835), .B2(n3672), .ZN(n2268)
         );
  OAI22_X2 U1792 ( .A1(n3475), .A2(n2837), .B1(n2836), .B2(n3673), .ZN(n2269)
         );
  OAI22_X2 U1793 ( .A1(n3474), .A2(n2838), .B1(n2837), .B2(n3672), .ZN(n2270)
         );
  OAI22_X2 U1794 ( .A1(n3474), .A2(n2839), .B1(n2838), .B2(n3672), .ZN(n2271)
         );
  OAI22_X2 U1795 ( .A1(n3475), .A2(n2840), .B1(n2839), .B2(n3672), .ZN(n2272)
         );
  OAI22_X2 U1796 ( .A1(n3474), .A2(n2841), .B1(n2840), .B2(n3672), .ZN(n2273)
         );
  OAI22_X2 U1797 ( .A1(n3474), .A2(n2842), .B1(n2841), .B2(n3673), .ZN(n2274)
         );
  OAI22_X2 U1798 ( .A1(n3475), .A2(n2843), .B1(n2842), .B2(n3673), .ZN(n2275)
         );
  OAI22_X2 U1799 ( .A1(n3474), .A2(n2844), .B1(n2843), .B2(n3672), .ZN(n2276)
         );
  OAI22_X2 U1800 ( .A1(n3474), .A2(n2845), .B1(n2844), .B2(n3673), .ZN(n2277)
         );
  OAI22_X2 U1803 ( .A1(n449), .A2(n2848), .B1(n2847), .B2(n3673), .ZN(n2280)
         );
  OAI22_X2 U1804 ( .A1(n449), .A2(n2849), .B1(n2848), .B2(n3672), .ZN(n2281)
         );
  OAI22_X2 U1805 ( .A1(n3474), .A2(n2850), .B1(n2849), .B2(n3673), .ZN(n2282)
         );
  OAI22_X2 U1806 ( .A1(n3475), .A2(n2851), .B1(n2850), .B2(n3673), .ZN(n2283)
         );
  OAI22_X2 U1808 ( .A1(n3475), .A2(n2853), .B1(n2852), .B2(n3672), .ZN(n2285)
         );
  OAI22_X2 U1809 ( .A1(n3475), .A2(n2854), .B1(n2853), .B2(n3673), .ZN(n2286)
         );
  OAI22_X2 U1810 ( .A1(n3474), .A2(n2855), .B1(n2854), .B2(n3672), .ZN(n2287)
         );
  OAI22_X2 U1811 ( .A1(n449), .A2(n2856), .B1(n2855), .B2(n3672), .ZN(n2288)
         );
  OAI22_X2 U1812 ( .A1(n3474), .A2(n2857), .B1(n2856), .B2(n3672), .ZN(n2289)
         );
  OAI22_X2 U1813 ( .A1(n3474), .A2(n2858), .B1(n2857), .B2(n3673), .ZN(n2290)
         );
  OAI22_X2 U1814 ( .A1(n3475), .A2(n2859), .B1(n2858), .B2(n3673), .ZN(n2291)
         );
  OAI22_X2 U1816 ( .A1(n3475), .A2(n2861), .B1(n2860), .B2(n3673), .ZN(n2293)
         );
  OAI22_X2 U1817 ( .A1(n3475), .A2(n2862), .B1(n2861), .B2(n3673), .ZN(n2294)
         );
  OAI22_X2 U1818 ( .A1(n3474), .A2(n2863), .B1(n2862), .B2(n3672), .ZN(n2295)
         );
  OAI22_X2 U1819 ( .A1(n3474), .A2(n2864), .B1(n2863), .B2(n3672), .ZN(n2296)
         );
  OAI22_X2 U1852 ( .A1(n446), .A2(n3283), .B1(n2898), .B2(n396), .ZN(n2067) );
  OAI22_X2 U1853 ( .A1(n446), .A2(n2866), .B1(n396), .B2(n3283), .ZN(n2299) );
  OAI22_X2 U1854 ( .A1(n3683), .A2(n2867), .B1(n2866), .B2(n396), .ZN(n2300)
         );
  OAI22_X2 U1855 ( .A1(n3683), .A2(n2868), .B1(n2867), .B2(n396), .ZN(n2301)
         );
  OAI22_X2 U1856 ( .A1(n446), .A2(n2869), .B1(n2868), .B2(n396), .ZN(n2302) );
  OAI22_X2 U1857 ( .A1(n3683), .A2(n2870), .B1(n2869), .B2(n396), .ZN(n2303)
         );
  OAI22_X2 U1858 ( .A1(n3683), .A2(n2871), .B1(n2870), .B2(n396), .ZN(n2304)
         );
  OAI22_X2 U1859 ( .A1(n446), .A2(n2872), .B1(n2871), .B2(n396), .ZN(n2305) );
  OAI22_X2 U1860 ( .A1(n3683), .A2(n2873), .B1(n2872), .B2(n396), .ZN(n2306)
         );
  OAI22_X2 U1861 ( .A1(n446), .A2(n2874), .B1(n2873), .B2(n396), .ZN(n2307) );
  OAI22_X2 U1862 ( .A1(n3683), .A2(n2875), .B1(n2874), .B2(n396), .ZN(n2308)
         );
  OAI22_X2 U1863 ( .A1(n3683), .A2(n2876), .B1(n2875), .B2(n396), .ZN(n2309)
         );
  OAI22_X2 U1865 ( .A1(n446), .A2(n2878), .B1(n2877), .B2(n396), .ZN(n2311) );
  OAI22_X2 U1866 ( .A1(n3683), .A2(n2879), .B1(n2878), .B2(n396), .ZN(n2312)
         );
  OAI22_X2 U1867 ( .A1(n3683), .A2(n2880), .B1(n2879), .B2(n396), .ZN(n2313)
         );
  OAI22_X2 U1868 ( .A1(n3683), .A2(n2881), .B1(n2880), .B2(n396), .ZN(n2314)
         );
  OAI22_X2 U1869 ( .A1(n446), .A2(n2882), .B1(n2881), .B2(n396), .ZN(n2315) );
  OAI22_X2 U1871 ( .A1(n3683), .A2(n2884), .B1(n2883), .B2(n396), .ZN(n2317)
         );
  OAI22_X2 U1872 ( .A1(n446), .A2(n2885), .B1(n2884), .B2(n396), .ZN(n2318) );
  OAI22_X2 U1873 ( .A1(n446), .A2(n2886), .B1(n2885), .B2(n396), .ZN(n2319) );
  OAI22_X2 U1874 ( .A1(n3683), .A2(n2887), .B1(n2886), .B2(n396), .ZN(n2320)
         );
  OAI22_X2 U1876 ( .A1(n446), .A2(n2889), .B1(n2888), .B2(n396), .ZN(n2322) );
  OAI22_X2 U1877 ( .A1(n3683), .A2(n2890), .B1(n2889), .B2(n396), .ZN(n2323)
         );
  OAI22_X2 U1878 ( .A1(n446), .A2(n2891), .B1(n2890), .B2(n396), .ZN(n2324) );
  OAI22_X2 U1879 ( .A1(n3683), .A2(n2892), .B1(n2891), .B2(n396), .ZN(n2325)
         );
  OAI22_X2 U1880 ( .A1(n446), .A2(n2893), .B1(n2892), .B2(n396), .ZN(n2326) );
  OAI22_X2 U1881 ( .A1(n446), .A2(n2894), .B1(n2893), .B2(n396), .ZN(n2327) );
  OAI22_X2 U1882 ( .A1(n446), .A2(n2895), .B1(n2894), .B2(n396), .ZN(n2328) );
  OAI22_X2 U1884 ( .A1(n3683), .A2(n2897), .B1(n2896), .B2(n396), .ZN(n2330)
         );
  OAI22_X2 U1982 ( .A1(n3459), .A2(n3689), .B1(n2964), .B2(n3698), .ZN(n2069)
         );
  OAI22_X2 U1983 ( .A1(n3459), .A2(n2932), .B1(n3698), .B2(n3689), .ZN(n2367)
         );
  OAI22_X2 U1984 ( .A1(n3459), .A2(n2933), .B1(n2932), .B2(n3698), .ZN(n2368)
         );
  OAI22_X2 U1985 ( .A1(n3459), .A2(n2934), .B1(n2933), .B2(n3698), .ZN(n2369)
         );
  OAI22_X2 U1986 ( .A1(n3459), .A2(n2935), .B1(n2934), .B2(n3698), .ZN(n2370)
         );
  OAI22_X2 U1987 ( .A1(n3459), .A2(n2936), .B1(n2935), .B2(n3698), .ZN(n2371)
         );
  OAI22_X2 U1988 ( .A1(n3459), .A2(n2937), .B1(n2936), .B2(n3698), .ZN(n2372)
         );
  OAI22_X2 U1989 ( .A1(n3459), .A2(n2938), .B1(n2937), .B2(n3698), .ZN(n2373)
         );
  OAI22_X2 U1990 ( .A1(n3458), .A2(n2939), .B1(n2938), .B2(n3698), .ZN(n2374)
         );
  OAI22_X2 U1991 ( .A1(n3459), .A2(n2940), .B1(n2939), .B2(n3698), .ZN(n2375)
         );
  OAI22_X2 U1992 ( .A1(n3459), .A2(n2941), .B1(n2940), .B2(n3698), .ZN(n2376)
         );
  OAI22_X2 U1993 ( .A1(n3458), .A2(n2942), .B1(n2941), .B2(n3698), .ZN(n2377)
         );
  OAI22_X2 U1994 ( .A1(n3459), .A2(n2943), .B1(n2942), .B2(n3698), .ZN(n2378)
         );
  OAI22_X2 U1995 ( .A1(n3459), .A2(n2944), .B1(n2943), .B2(n3698), .ZN(n2379)
         );
  OAI22_X2 U1996 ( .A1(n3459), .A2(n2945), .B1(n2944), .B2(n3698), .ZN(n2380)
         );
  OAI22_X2 U1997 ( .A1(n3459), .A2(n2946), .B1(n2945), .B2(n3698), .ZN(n2381)
         );
  OAI22_X2 U1998 ( .A1(n3458), .A2(n2947), .B1(n2946), .B2(n3698), .ZN(n2382)
         );
  OAI22_X2 U1999 ( .A1(n3458), .A2(n2948), .B1(n2947), .B2(n3698), .ZN(n2383)
         );
  OAI22_X2 U2001 ( .A1(n3459), .A2(n2950), .B1(n2949), .B2(n3698), .ZN(n2385)
         );
  OAI22_X2 U2002 ( .A1(n3459), .A2(n2951), .B1(n2950), .B2(n3698), .ZN(n2386)
         );
  OAI22_X2 U2003 ( .A1(n3459), .A2(n2952), .B1(n2951), .B2(n3698), .ZN(n2387)
         );
  OAI22_X2 U2004 ( .A1(n3459), .A2(n2953), .B1(n2952), .B2(n3698), .ZN(n2388)
         );
  OAI22_X2 U2006 ( .A1(n3459), .A2(n2955), .B1(n2954), .B2(n3698), .ZN(n2390)
         );
  OAI22_X2 U2007 ( .A1(n3459), .A2(n2956), .B1(n2955), .B2(n3698), .ZN(n2391)
         );
  OAI22_X2 U2008 ( .A1(n3459), .A2(n2957), .B1(n2956), .B2(n3698), .ZN(n2392)
         );
  OAI22_X2 U2009 ( .A1(n3459), .A2(n2958), .B1(n2957), .B2(n3698), .ZN(n2393)
         );
  OAI22_X2 U2010 ( .A1(n3459), .A2(n2959), .B1(n2958), .B2(n3698), .ZN(n2394)
         );
  OAI22_X2 U2011 ( .A1(n3459), .A2(n2960), .B1(n2959), .B2(n3698), .ZN(n2395)
         );
  OAI22_X2 U2012 ( .A1(n3459), .A2(n2961), .B1(n2960), .B2(n3698), .ZN(n2396)
         );
  OAI22_X2 U2013 ( .A1(n3459), .A2(n2962), .B1(n2961), .B2(n3698), .ZN(n2397)
         );
  OAI22_X2 U2014 ( .A1(n3459), .A2(n2963), .B1(n2962), .B2(n3698), .ZN(n2398)
         );
  OAI22_X2 U2047 ( .A1(n3667), .A2(n3286), .B1(n2997), .B2(n3571), .ZN(n2070)
         );
  OAI22_X2 U2049 ( .A1(n3667), .A2(n2966), .B1(n2965), .B2(n3571), .ZN(n2402)
         );
  OAI22_X2 U2052 ( .A1(n3667), .A2(n2969), .B1(n2968), .B2(n3571), .ZN(n2405)
         );
  OAI22_X2 U2054 ( .A1(n3667), .A2(n2971), .B1(n2970), .B2(n3571), .ZN(n2407)
         );
  OAI22_X2 U2057 ( .A1(n3667), .A2(n2974), .B1(n2973), .B2(n3571), .ZN(n2410)
         );
  OAI22_X2 U2065 ( .A1(n3667), .A2(n2982), .B1(n2981), .B2(n3571), .ZN(n2418)
         );
  OAI22_X2 U2069 ( .A1(n3667), .A2(n2986), .B1(n2985), .B2(n3571), .ZN(n2422)
         );
  OAI22_X2 U2072 ( .A1(n3667), .A2(n2989), .B1(n2988), .B2(n3571), .ZN(n2425)
         );
  OAI22_X2 U2073 ( .A1(n3667), .A2(n2990), .B1(n2989), .B2(n3571), .ZN(n2426)
         );
  OAI22_X2 U2074 ( .A1(n3667), .A2(n2991), .B1(n2990), .B2(n3571), .ZN(n2427)
         );
  OAI22_X2 U2076 ( .A1(n3667), .A2(n2993), .B1(n2992), .B2(n3571), .ZN(n2429)
         );
  OAI22_X2 U2077 ( .A1(n3667), .A2(n2994), .B1(n2993), .B2(n3571), .ZN(n2430)
         );
  OAI22_X2 U2078 ( .A1(n3667), .A2(n2995), .B1(n2994), .B2(n3571), .ZN(n2431)
         );
  OAI22_X2 U2079 ( .A1(n3667), .A2(n2996), .B1(n2995), .B2(n3571), .ZN(n2432)
         );
  OAI22_X2 U2124 ( .A1(n3552), .A2(n3009), .B1(n3008), .B2(n3567), .ZN(n2446)
         );
  OAI22_X2 U2179 ( .A1(n431), .A2(n3032), .B1(n3031), .B2(n381), .ZN(n2470) );
  OAI22_X2 U2183 ( .A1(n431), .A2(n3036), .B1(n3035), .B2(n381), .ZN(n2474) );
  OAI22_X2 U2184 ( .A1(n431), .A2(n3037), .B1(n3036), .B2(n381), .ZN(n2475) );
  OAI22_X2 U2188 ( .A1(n431), .A2(n3041), .B1(n381), .B2(n3040), .ZN(n2479) );
  OAI22_X2 U2190 ( .A1(n431), .A2(n3043), .B1(n3042), .B2(n381), .ZN(n2481) );
  OAI22_X2 U2197 ( .A1(n431), .A2(n3050), .B1(n3049), .B2(n381), .ZN(n2488) );
  OAI22_X2 U2202 ( .A1(n431), .A2(n3055), .B1(n3054), .B2(n381), .ZN(n2493) );
  OAI22_X2 U2205 ( .A1(n431), .A2(n3058), .B1(n3057), .B2(n381), .ZN(n2496) );
  OAI22_X2 U2207 ( .A1(n431), .A2(n3060), .B1(n3059), .B2(n381), .ZN(n2498) );
  OAI22_X2 U2242 ( .A1(n428), .A2(n3289), .B1(n3096), .B2(n3664), .ZN(n2073)
         );
  OAI22_X2 U2247 ( .A1(n428), .A2(n3068), .B1(n3067), .B2(n3664), .ZN(n2507)
         );
  OAI22_X2 U2248 ( .A1(n428), .A2(n3069), .B1(n3068), .B2(n3664), .ZN(n2508)
         );
  OAI22_X2 U2249 ( .A1(n428), .A2(n3070), .B1(n3069), .B2(n3664), .ZN(n2509)
         );
  OAI22_X2 U2250 ( .A1(n428), .A2(n3071), .B1(n3070), .B2(n3664), .ZN(n2510)
         );
  OAI22_X2 U2251 ( .A1(n428), .A2(n3072), .B1(n3071), .B2(n3664), .ZN(n2511)
         );
  OAI22_X2 U2252 ( .A1(n428), .A2(n3073), .B1(n3072), .B2(n3664), .ZN(n2512)
         );
  OAI22_X2 U2253 ( .A1(n428), .A2(n3074), .B1(n3073), .B2(n3664), .ZN(n2513)
         );
  OAI22_X2 U2254 ( .A1(n428), .A2(n3075), .B1(n3074), .B2(n3664), .ZN(n2514)
         );
  OAI22_X2 U2255 ( .A1(n428), .A2(n3076), .B1(n3075), .B2(n3664), .ZN(n2515)
         );
  OAI22_X2 U2256 ( .A1(n428), .A2(n3077), .B1(n3076), .B2(n3664), .ZN(n2516)
         );
  OAI22_X2 U2257 ( .A1(n428), .A2(n3078), .B1(n3077), .B2(n3664), .ZN(n2517)
         );
  OAI22_X2 U2258 ( .A1(n428), .A2(n3079), .B1(n3078), .B2(n3664), .ZN(n2518)
         );
  OAI22_X2 U2260 ( .A1(n428), .A2(n3081), .B1(n3080), .B2(n3664), .ZN(n2520)
         );
  OAI22_X2 U2261 ( .A1(n428), .A2(n3082), .B1(n3081), .B2(n3664), .ZN(n2521)
         );
  OAI22_X2 U2262 ( .A1(n428), .A2(n3083), .B1(n3082), .B2(n3664), .ZN(n2522)
         );
  OAI22_X2 U2263 ( .A1(n428), .A2(n3084), .B1(n3083), .B2(n3664), .ZN(n2523)
         );
  OAI22_X2 U2264 ( .A1(n428), .A2(n3085), .B1(n3084), .B2(n3664), .ZN(n2524)
         );
  OAI22_X2 U2265 ( .A1(n428), .A2(n3086), .B1(n3085), .B2(n3664), .ZN(n2525)
         );
  OAI22_X2 U2267 ( .A1(n428), .A2(n3088), .B1(n3087), .B2(n3664), .ZN(n2527)
         );
  OAI22_X2 U2268 ( .A1(n428), .A2(n3089), .B1(n3088), .B2(n3664), .ZN(n2528)
         );
  OAI22_X2 U2269 ( .A1(n428), .A2(n3090), .B1(n3089), .B2(n3664), .ZN(n2529)
         );
  OAI22_X2 U2270 ( .A1(n428), .A2(n3091), .B1(n3090), .B2(n3664), .ZN(n2530)
         );
  OAI22_X2 U2271 ( .A1(n428), .A2(n3092), .B1(n3091), .B2(n3664), .ZN(n2531)
         );
  OAI22_X2 U2272 ( .A1(n428), .A2(n3093), .B1(n3092), .B2(n3664), .ZN(n2532)
         );
  OAI22_X2 U2273 ( .A1(n428), .A2(n3094), .B1(n3093), .B2(n3664), .ZN(n2533)
         );
  OAI22_X2 U2274 ( .A1(n428), .A2(n3095), .B1(n3094), .B2(n3664), .ZN(n2534)
         );
  OAI22_X2 U2308 ( .A1(n425), .A2(n3097), .B1(n3533), .B2(n3290), .ZN(n2537)
         );
  OAI22_X2 U2309 ( .A1(n425), .A2(n3098), .B1(n3097), .B2(n3533), .ZN(n2538)
         );
  OAI22_X2 U2375 ( .A1(n422), .A2(n3132), .B1(n3131), .B2(n372), .ZN(n2573) );
  OAI22_X2 U2377 ( .A1(n422), .A2(n3134), .B1(n3133), .B2(n372), .ZN(n2575) );
  OAI22_X2 U2378 ( .A1(n422), .A2(n3135), .B1(n3134), .B2(n372), .ZN(n2576) );
  OAI22_X2 U2379 ( .A1(n422), .A2(n3136), .B1(n3135), .B2(n372), .ZN(n2577) );
  OAI22_X2 U2382 ( .A1(n422), .A2(n3139), .B1(n3138), .B2(n372), .ZN(n2580) );
  OAI22_X2 U2383 ( .A1(n422), .A2(n3140), .B1(n3139), .B2(n372), .ZN(n2581) );
  OAI22_X2 U2384 ( .A1(n422), .A2(n3141), .B1(n3140), .B2(n372), .ZN(n2582) );
  OAI22_X2 U2386 ( .A1(n422), .A2(n3143), .B1(n3142), .B2(n372), .ZN(n2584) );
  OAI22_X2 U2387 ( .A1(n422), .A2(n3144), .B1(n3143), .B2(n372), .ZN(n2585) );
  OAI22_X2 U2388 ( .A1(n422), .A2(n3145), .B1(n3144), .B2(n372), .ZN(n2586) );
  OAI22_X2 U2389 ( .A1(n422), .A2(n3146), .B1(n3145), .B2(n372), .ZN(n2587) );
  OAI22_X2 U2392 ( .A1(n422), .A2(n3149), .B1(n3148), .B2(n372), .ZN(n2590) );
  OAI22_X2 U2393 ( .A1(n422), .A2(n3150), .B1(n3149), .B2(n372), .ZN(n2591) );
  OAI22_X2 U2437 ( .A1(n3526), .A2(n3292), .B1(n3195), .B2(n3511), .ZN(n2076)
         );
  OAI22_X2 U2461 ( .A1(n3526), .A2(n3186), .B1(n3185), .B2(n3511), .ZN(n2628)
         );
  OAI22_X2 U2465 ( .A1(n3526), .A2(n3190), .B1(n3189), .B2(n3511), .ZN(n2632)
         );
  OAI22_X2 U2466 ( .A1(n3526), .A2(n3191), .B1(n3190), .B2(n3511), .ZN(n2633)
         );
  OAI22_X2 U2467 ( .A1(n3526), .A2(n3192), .B1(n3191), .B2(n3511), .ZN(n2634)
         );
  OAI22_X2 U2468 ( .A1(n3526), .A2(n3193), .B1(n3192), .B2(n3511), .ZN(n2635)
         );
  OAI22_X2 U2469 ( .A1(n3526), .A2(n3194), .B1(n3193), .B2(n3511), .ZN(n2636)
         );
  NAND2_X4 U2568 ( .A1(n3239), .A2(n381), .ZN(n431) );
  XOR2_X2 U2569 ( .A(a[8]), .B(n333), .Z(n3239) );
  NAND2_X1 U2585 ( .A1(n3749), .A2(n324), .ZN(n3677) );
  XNOR2_X1 U2586 ( .A(n3741), .B(n351), .ZN(n3588) );
  INV_X4 U2587 ( .A(a[20]), .ZN(n3741) );
  INV_X2 U2588 ( .A(n3553), .ZN(n3554) );
  INV_X2 U2589 ( .A(n3573), .ZN(n3574) );
  INV_X1 U2590 ( .A(n336), .ZN(n3668) );
  INV_X1 U2591 ( .A(n357), .ZN(n3730) );
  INV_X1 U2592 ( .A(n366), .ZN(n416) );
  INV_X1 U2593 ( .A(n330), .ZN(n3289) );
  INV_X1 U2594 ( .A(n330), .ZN(n3659) );
  INV_X1 U2595 ( .A(n321), .ZN(n3292) );
  INV_X1 U2596 ( .A(n321), .ZN(n3597) );
  INV_X1 U2597 ( .A(n354), .ZN(n3281) );
  INV_X1 U2598 ( .A(n354), .ZN(n3633) );
  INV_X4 U2599 ( .A(a[30]), .ZN(n3745) );
  INV_X2 U2600 ( .A(a[6]), .ZN(n3737) );
  INV_X4 U2601 ( .A(a[4]), .ZN(n3749) );
  INV_X2 U2602 ( .A(a[26]), .ZN(n3657) );
  INV_X4 U2603 ( .A(a[22]), .ZN(n3614) );
  INV_X2 U2604 ( .A(a[28]), .ZN(n3604) );
  XOR2_X1 U2605 ( .A(a[28]), .B(n363), .Z(n3229) );
  INV_X4 U2606 ( .A(a[24]), .ZN(n3472) );
  XOR2_X1 U2607 ( .A(a[10]), .B(n336), .Z(n3238) );
  INV_X2 U2608 ( .A(a[10]), .ZN(n3624) );
  INV_X1 U2609 ( .A(a[16]), .ZN(n3688) );
  NAND2_X1 U2610 ( .A1(a[2]), .A2(n321), .ZN(n3598) );
  INV_X2 U2611 ( .A(a[0]), .ZN(n369) );
  INV_X1 U2612 ( .A(n360), .ZN(n3573) );
  NAND2_X1 U2613 ( .A1(n3604), .A2(n360), .ZN(n3606) );
  XOR2_X1 U2614 ( .A(a[26]), .B(n360), .Z(n3230) );
  INV_X1 U2615 ( .A(n529), .ZN(n2637) );
  XNOR2_X1 U2616 ( .A(n529), .B(n366), .ZN(n2668) );
  XNOR2_X1 U2617 ( .A(n529), .B(n363), .ZN(n2701) );
  XNOR2_X1 U2618 ( .A(n529), .B(n3574), .ZN(n2734) );
  XNOR2_X1 U2619 ( .A(n529), .B(n3731), .ZN(n2767) );
  XNOR2_X1 U2620 ( .A(n529), .B(n348), .ZN(n2866) );
  XNOR2_X1 U2621 ( .A(n529), .B(n324), .ZN(n3130) );
  XNOR2_X1 U2622 ( .A(n529), .B(n336), .ZN(n2998) );
  XNOR2_X1 U2623 ( .A(n529), .B(n354), .ZN(n2800) );
  XNOR2_X1 U2624 ( .A(n529), .B(n345), .ZN(n2899) );
  XNOR2_X1 U2625 ( .A(n529), .B(n3554), .ZN(n3031) );
  XNOR2_X1 U2626 ( .A(n529), .B(n342), .ZN(n2932) );
  XNOR2_X1 U2627 ( .A(n529), .B(n351), .ZN(n2833) );
  XNOR2_X1 U2628 ( .A(n529), .B(n339), .ZN(n2965) );
  XNOR2_X1 U2629 ( .A(n529), .B(n330), .ZN(n3064) );
  XNOR2_X1 U2630 ( .A(n529), .B(n321), .ZN(n3163) );
  XNOR2_X1 U2631 ( .A(n529), .B(n327), .ZN(n3097) );
  INV_X1 U2632 ( .A(n527), .ZN(n2638) );
  XNOR2_X1 U2633 ( .A(n527), .B(n366), .ZN(n2669) );
  XNOR2_X1 U2634 ( .A(n527), .B(n363), .ZN(n2702) );
  XNOR2_X1 U2635 ( .A(n527), .B(n3574), .ZN(n2735) );
  XNOR2_X1 U2636 ( .A(n527), .B(n3669), .ZN(n2999) );
  XNOR2_X1 U2637 ( .A(n527), .B(n357), .ZN(n2768) );
  XNOR2_X1 U2638 ( .A(n527), .B(n351), .ZN(n2834) );
  XNOR2_X1 U2639 ( .A(n527), .B(n324), .ZN(n3131) );
  XNOR2_X1 U2640 ( .A(n527), .B(n354), .ZN(n2801) );
  XNOR2_X1 U2641 ( .A(n527), .B(n345), .ZN(n2900) );
  XNOR2_X1 U2642 ( .A(n527), .B(n339), .ZN(n2966) );
  XNOR2_X1 U2643 ( .A(n527), .B(n348), .ZN(n2867) );
  XNOR2_X1 U2644 ( .A(n527), .B(n342), .ZN(n2933) );
  XNOR2_X1 U2645 ( .A(n527), .B(n327), .ZN(n3098) );
  XNOR2_X1 U2646 ( .A(n527), .B(n330), .ZN(n3065) );
  XNOR2_X1 U2647 ( .A(n527), .B(n321), .ZN(n3164) );
  INV_X1 U2648 ( .A(n525), .ZN(n2639) );
  XNOR2_X1 U2649 ( .A(n525), .B(n366), .ZN(n2670) );
  XNOR2_X1 U2650 ( .A(n525), .B(n363), .ZN(n2703) );
  XNOR2_X1 U2651 ( .A(n525), .B(n3574), .ZN(n2736) );
  XNOR2_X1 U2652 ( .A(n525), .B(n351), .ZN(n2835) );
  XNOR2_X1 U2653 ( .A(n525), .B(n336), .ZN(n3000) );
  XNOR2_X1 U2654 ( .A(n525), .B(n339), .ZN(n2967) );
  XNOR2_X1 U2655 ( .A(n525), .B(n354), .ZN(n2802) );
  XNOR2_X1 U2656 ( .A(n525), .B(n345), .ZN(n2901) );
  XNOR2_X1 U2657 ( .A(n525), .B(n342), .ZN(n2934) );
  XNOR2_X1 U2658 ( .A(n525), .B(n357), .ZN(n2769) );
  XNOR2_X1 U2659 ( .A(n525), .B(n348), .ZN(n2868) );
  XNOR2_X1 U2660 ( .A(n525), .B(n327), .ZN(n3099) );
  XNOR2_X1 U2661 ( .A(n525), .B(n330), .ZN(n3066) );
  XNOR2_X1 U2662 ( .A(n525), .B(n321), .ZN(n3165) );
  XNOR2_X1 U2663 ( .A(n525), .B(n324), .ZN(n3132) );
  INV_X1 U2664 ( .A(n523), .ZN(n2640) );
  XNOR2_X1 U2665 ( .A(n523), .B(n366), .ZN(n2671) );
  XNOR2_X1 U2666 ( .A(n523), .B(n363), .ZN(n2704) );
  XNOR2_X1 U2667 ( .A(n523), .B(n3574), .ZN(n2737) );
  XNOR2_X1 U2668 ( .A(n523), .B(n354), .ZN(n2803) );
  XNOR2_X1 U2669 ( .A(n523), .B(n3647), .ZN(n2968) );
  XNOR2_X1 U2670 ( .A(n523), .B(n342), .ZN(n2935) );
  XNOR2_X1 U2671 ( .A(n523), .B(n327), .ZN(n3100) );
  XNOR2_X1 U2672 ( .A(n523), .B(n321), .ZN(n3166) );
  XNOR2_X1 U2673 ( .A(n523), .B(n357), .ZN(n2770) );
  XNOR2_X1 U2674 ( .A(n523), .B(n348), .ZN(n2869) );
  XNOR2_X1 U2675 ( .A(n523), .B(n345), .ZN(n2902) );
  XNOR2_X1 U2676 ( .A(n523), .B(n330), .ZN(n3067) );
  XNOR2_X1 U2677 ( .A(n523), .B(n351), .ZN(n2836) );
  XNOR2_X1 U2678 ( .A(n523), .B(n324), .ZN(n3133) );
  XNOR2_X1 U2679 ( .A(n523), .B(n3554), .ZN(n3034) );
  INV_X1 U2680 ( .A(n521), .ZN(n2641) );
  XNOR2_X1 U2681 ( .A(n521), .B(n366), .ZN(n2672) );
  XNOR2_X1 U2682 ( .A(n521), .B(n363), .ZN(n2705) );
  XNOR2_X1 U2683 ( .A(n521), .B(n342), .ZN(n2936) );
  XNOR2_X1 U2684 ( .A(n521), .B(n357), .ZN(n2771) );
  XNOR2_X1 U2685 ( .A(n521), .B(n321), .ZN(n3167) );
  XNOR2_X1 U2686 ( .A(n521), .B(n345), .ZN(n2903) );
  XNOR2_X1 U2687 ( .A(n521), .B(n354), .ZN(n2804) );
  XNOR2_X1 U2688 ( .A(n521), .B(n327), .ZN(n3101) );
  XNOR2_X1 U2689 ( .A(n521), .B(n348), .ZN(n2870) );
  XNOR2_X1 U2690 ( .A(n521), .B(n3574), .ZN(n2738) );
  XNOR2_X1 U2691 ( .A(n521), .B(n351), .ZN(n2837) );
  XNOR2_X1 U2692 ( .A(n521), .B(n330), .ZN(n3068) );
  XNOR2_X1 U2693 ( .A(n521), .B(n324), .ZN(n3134) );
  XNOR2_X1 U2694 ( .A(n521), .B(n3554), .ZN(n3035) );
  XNOR2_X1 U2695 ( .A(n521), .B(n339), .ZN(n2969) );
  INV_X1 U2696 ( .A(n519), .ZN(n2642) );
  XNOR2_X1 U2697 ( .A(n519), .B(n366), .ZN(n2673) );
  XNOR2_X1 U2698 ( .A(n519), .B(n363), .ZN(n2706) );
  XNOR2_X1 U2699 ( .A(n519), .B(n342), .ZN(n2937) );
  XNOR2_X1 U2700 ( .A(n519), .B(n345), .ZN(n2904) );
  XNOR2_X1 U2701 ( .A(n519), .B(n357), .ZN(n2772) );
  XNOR2_X1 U2702 ( .A(n519), .B(n330), .ZN(n3069) );
  XNOR2_X1 U2703 ( .A(n519), .B(n336), .ZN(n3003) );
  XNOR2_X1 U2704 ( .A(n519), .B(n321), .ZN(n3168) );
  XNOR2_X1 U2705 ( .A(n519), .B(n3574), .ZN(n2739) );
  XNOR2_X1 U2706 ( .A(n519), .B(n3554), .ZN(n3036) );
  XNOR2_X1 U2707 ( .A(n519), .B(n354), .ZN(n2805) );
  XNOR2_X1 U2708 ( .A(n519), .B(n351), .ZN(n2838) );
  XNOR2_X1 U2709 ( .A(n519), .B(n348), .ZN(n2871) );
  XNOR2_X1 U2710 ( .A(n519), .B(n327), .ZN(n3102) );
  XNOR2_X1 U2711 ( .A(n519), .B(n339), .ZN(n2970) );
  XNOR2_X1 U2712 ( .A(n519), .B(n324), .ZN(n3135) );
  INV_X1 U2713 ( .A(n515), .ZN(n2644) );
  XNOR2_X1 U2714 ( .A(n515), .B(n363), .ZN(n2708) );
  XNOR2_X1 U2715 ( .A(n515), .B(n366), .ZN(n2675) );
  XNOR2_X1 U2716 ( .A(n515), .B(n345), .ZN(n2906) );
  XNOR2_X1 U2717 ( .A(n515), .B(n3731), .ZN(n2774) );
  XNOR2_X1 U2718 ( .A(n515), .B(n3574), .ZN(n2741) );
  XNOR2_X1 U2719 ( .A(n515), .B(n348), .ZN(n2873) );
  XNOR2_X1 U2720 ( .A(n515), .B(n324), .ZN(n3137) );
  XNOR2_X1 U2721 ( .A(n515), .B(n351), .ZN(n2840) );
  XNOR2_X1 U2722 ( .A(n515), .B(n327), .ZN(n3104) );
  XNOR2_X1 U2723 ( .A(n515), .B(n354), .ZN(n2807) );
  XNOR2_X1 U2724 ( .A(n515), .B(n3554), .ZN(n3038) );
  XNOR2_X1 U2725 ( .A(n515), .B(n330), .ZN(n3071) );
  XNOR2_X1 U2726 ( .A(n515), .B(n342), .ZN(n2939) );
  XNOR2_X1 U2727 ( .A(n515), .B(n321), .ZN(n3170) );
  XNOR2_X1 U2728 ( .A(n515), .B(n336), .ZN(n3005) );
  XNOR2_X1 U2729 ( .A(n515), .B(n339), .ZN(n2972) );
  INV_X1 U2730 ( .A(n517), .ZN(n2643) );
  XNOR2_X1 U2731 ( .A(n517), .B(n366), .ZN(n2674) );
  XNOR2_X1 U2732 ( .A(n517), .B(n363), .ZN(n2707) );
  XNOR2_X1 U2733 ( .A(n517), .B(n3731), .ZN(n2773) );
  XNOR2_X1 U2734 ( .A(n517), .B(n345), .ZN(n2905) );
  XNOR2_X1 U2735 ( .A(n517), .B(n348), .ZN(n2872) );
  XNOR2_X1 U2736 ( .A(n517), .B(n3574), .ZN(n2740) );
  XNOR2_X1 U2737 ( .A(n517), .B(n3554), .ZN(n3037) );
  XNOR2_X1 U2738 ( .A(n517), .B(n330), .ZN(n3070) );
  XNOR2_X1 U2739 ( .A(n517), .B(n351), .ZN(n2839) );
  XNOR2_X1 U2740 ( .A(n517), .B(n324), .ZN(n3136) );
  XNOR2_X1 U2741 ( .A(n517), .B(n336), .ZN(n3004) );
  XNOR2_X1 U2742 ( .A(n517), .B(n327), .ZN(n3103) );
  XNOR2_X1 U2743 ( .A(n517), .B(n354), .ZN(n2806) );
  XNOR2_X1 U2744 ( .A(n517), .B(n342), .ZN(n2938) );
  XNOR2_X1 U2745 ( .A(n517), .B(n321), .ZN(n3169) );
  XNOR2_X1 U2746 ( .A(n517), .B(n339), .ZN(n2971) );
  INV_X1 U2747 ( .A(n513), .ZN(n2645) );
  XNOR2_X1 U2748 ( .A(n513), .B(n3574), .ZN(n2742) );
  XNOR2_X1 U2749 ( .A(n513), .B(n363), .ZN(n2709) );
  XNOR2_X1 U2750 ( .A(n513), .B(n348), .ZN(n2874) );
  XNOR2_X1 U2751 ( .A(n513), .B(n357), .ZN(n2775) );
  XNOR2_X1 U2752 ( .A(n513), .B(n342), .ZN(n2940) );
  XNOR2_X1 U2753 ( .A(n513), .B(n354), .ZN(n2808) );
  XNOR2_X1 U2754 ( .A(n513), .B(n339), .ZN(n2973) );
  XNOR2_X1 U2755 ( .A(n513), .B(n351), .ZN(n2841) );
  XNOR2_X1 U2756 ( .A(n513), .B(n3554), .ZN(n3039) );
  XNOR2_X1 U2757 ( .A(n513), .B(n324), .ZN(n3138) );
  XNOR2_X1 U2758 ( .A(n513), .B(n366), .ZN(n2676) );
  XNOR2_X1 U2759 ( .A(n513), .B(n321), .ZN(n3171) );
  XNOR2_X1 U2760 ( .A(n513), .B(n330), .ZN(n3072) );
  XNOR2_X1 U2761 ( .A(n513), .B(n336), .ZN(n3006) );
  XNOR2_X1 U2762 ( .A(n513), .B(n345), .ZN(n2907) );
  XNOR2_X1 U2763 ( .A(n513), .B(n327), .ZN(n3105) );
  INV_X1 U2764 ( .A(n511), .ZN(n2646) );
  XNOR2_X1 U2765 ( .A(n511), .B(n3574), .ZN(n2743) );
  XNOR2_X1 U2766 ( .A(n511), .B(n363), .ZN(n2710) );
  XNOR2_X1 U2767 ( .A(n511), .B(n348), .ZN(n2875) );
  XNOR2_X1 U2768 ( .A(n511), .B(n336), .ZN(n3007) );
  XNOR2_X1 U2769 ( .A(n511), .B(n339), .ZN(n2974) );
  XNOR2_X1 U2770 ( .A(n511), .B(n357), .ZN(n2776) );
  XNOR2_X1 U2771 ( .A(n511), .B(n321), .ZN(n3172) );
  XNOR2_X1 U2772 ( .A(n511), .B(n366), .ZN(n2677) );
  XNOR2_X1 U2773 ( .A(n511), .B(n351), .ZN(n2842) );
  XNOR2_X1 U2774 ( .A(n511), .B(n330), .ZN(n3073) );
  XNOR2_X1 U2775 ( .A(n511), .B(n324), .ZN(n3139) );
  XNOR2_X1 U2776 ( .A(n511), .B(n327), .ZN(n3106) );
  XNOR2_X1 U2777 ( .A(n511), .B(n345), .ZN(n2908) );
  XNOR2_X1 U2778 ( .A(n511), .B(n342), .ZN(n2941) );
  XNOR2_X1 U2779 ( .A(n511), .B(n354), .ZN(n2809) );
  INV_X1 U2780 ( .A(n507), .ZN(n2648) );
  XNOR2_X1 U2781 ( .A(n507), .B(n363), .ZN(n2712) );
  XNOR2_X1 U2782 ( .A(n507), .B(n366), .ZN(n2679) );
  XNOR2_X1 U2783 ( .A(n507), .B(n3574), .ZN(n2745) );
  XNOR2_X1 U2784 ( .A(n507), .B(n339), .ZN(n2976) );
  XNOR2_X1 U2785 ( .A(n507), .B(n330), .ZN(n3075) );
  XNOR2_X1 U2786 ( .A(n507), .B(n336), .ZN(n3009) );
  XNOR2_X1 U2787 ( .A(n507), .B(n324), .ZN(n3141) );
  XNOR2_X1 U2788 ( .A(n507), .B(n354), .ZN(n2811) );
  XNOR2_X1 U2789 ( .A(n507), .B(n348), .ZN(n2877) );
  XNOR2_X1 U2790 ( .A(n507), .B(n321), .ZN(n3174) );
  XNOR2_X1 U2791 ( .A(n507), .B(n342), .ZN(n2943) );
  XNOR2_X1 U2792 ( .A(n507), .B(n327), .ZN(n3108) );
  XNOR2_X1 U2793 ( .A(n507), .B(n357), .ZN(n2778) );
  XNOR2_X1 U2794 ( .A(n507), .B(n351), .ZN(n2844) );
  XNOR2_X1 U2795 ( .A(n507), .B(n345), .ZN(n2910) );
  INV_X1 U2796 ( .A(n509), .ZN(n2647) );
  XNOR2_X1 U2797 ( .A(n509), .B(n363), .ZN(n2711) );
  XNOR2_X1 U2798 ( .A(n509), .B(n3574), .ZN(n2744) );
  XNOR2_X1 U2799 ( .A(n509), .B(n366), .ZN(n2678) );
  XNOR2_X1 U2800 ( .A(n509), .B(n321), .ZN(n3173) );
  XNOR2_X1 U2801 ( .A(n509), .B(n336), .ZN(n3008) );
  XNOR2_X1 U2802 ( .A(n509), .B(n330), .ZN(n3074) );
  XNOR2_X1 U2803 ( .A(n509), .B(n351), .ZN(n2843) );
  XNOR2_X1 U2804 ( .A(n509), .B(n357), .ZN(n2777) );
  XNOR2_X1 U2805 ( .A(n509), .B(n339), .ZN(n2975) );
  XNOR2_X1 U2806 ( .A(n509), .B(n327), .ZN(n3107) );
  XNOR2_X1 U2807 ( .A(n509), .B(n324), .ZN(n3140) );
  XNOR2_X1 U2808 ( .A(n509), .B(n345), .ZN(n2909) );
  XNOR2_X1 U2809 ( .A(n509), .B(n348), .ZN(n2876) );
  XNOR2_X1 U2810 ( .A(n509), .B(n354), .ZN(n2810) );
  XNOR2_X1 U2811 ( .A(n509), .B(n3554), .ZN(n3041) );
  XNOR2_X1 U2812 ( .A(n509), .B(n342), .ZN(n2942) );
  INV_X1 U2813 ( .A(n505), .ZN(n2649) );
  XNOR2_X1 U2814 ( .A(n505), .B(n3669), .ZN(n3010) );
  XNOR2_X1 U2815 ( .A(n505), .B(n366), .ZN(n2680) );
  XNOR2_X1 U2816 ( .A(n505), .B(n363), .ZN(n2713) );
  XNOR2_X1 U2817 ( .A(n505), .B(n324), .ZN(n3142) );
  XNOR2_X1 U2818 ( .A(n505), .B(n354), .ZN(n2812) );
  XNOR2_X1 U2819 ( .A(n505), .B(n342), .ZN(n2944) );
  XNOR2_X1 U2820 ( .A(n505), .B(n3574), .ZN(n2746) );
  XNOR2_X1 U2821 ( .A(n505), .B(n321), .ZN(n3175) );
  XNOR2_X1 U2822 ( .A(n505), .B(n327), .ZN(n3109) );
  XNOR2_X1 U2823 ( .A(n505), .B(n357), .ZN(n2779) );
  XNOR2_X1 U2824 ( .A(n505), .B(n351), .ZN(n2845) );
  XNOR2_X1 U2825 ( .A(n505), .B(n348), .ZN(n2878) );
  XNOR2_X1 U2826 ( .A(n505), .B(n339), .ZN(n2977) );
  XNOR2_X1 U2827 ( .A(n505), .B(n330), .ZN(n3076) );
  XNOR2_X1 U2828 ( .A(n505), .B(n345), .ZN(n2911) );
  XNOR2_X1 U2829 ( .A(n505), .B(n3554), .ZN(n3043) );
  INV_X1 U2830 ( .A(n503), .ZN(n2650) );
  XNOR2_X1 U2831 ( .A(n503), .B(n363), .ZN(n2714) );
  XNOR2_X1 U2832 ( .A(n503), .B(n354), .ZN(n2813) );
  XNOR2_X1 U2833 ( .A(n503), .B(n327), .ZN(n3110) );
  XNOR2_X1 U2834 ( .A(n503), .B(n342), .ZN(n2945) );
  XNOR2_X1 U2835 ( .A(n503), .B(n366), .ZN(n2681) );
  XNOR2_X1 U2836 ( .A(n503), .B(n321), .ZN(n3176) );
  XNOR2_X1 U2837 ( .A(n503), .B(n324), .ZN(n3143) );
  XNOR2_X1 U2838 ( .A(n503), .B(n351), .ZN(n2846) );
  XNOR2_X1 U2839 ( .A(n503), .B(n345), .ZN(n2912) );
  XNOR2_X1 U2840 ( .A(n503), .B(n357), .ZN(n2780) );
  XNOR2_X1 U2841 ( .A(n503), .B(n3554), .ZN(n3044) );
  XNOR2_X1 U2842 ( .A(n503), .B(n336), .ZN(n3011) );
  XNOR2_X1 U2843 ( .A(n503), .B(n330), .ZN(n3077) );
  XNOR2_X1 U2844 ( .A(n503), .B(n3574), .ZN(n2747) );
  XNOR2_X1 U2845 ( .A(n503), .B(n348), .ZN(n2879) );
  XNOR2_X1 U2846 ( .A(n503), .B(n339), .ZN(n2978) );
  INV_X1 U2847 ( .A(n499), .ZN(n2652) );
  XNOR2_X1 U2848 ( .A(n499), .B(n357), .ZN(n2782) );
  XNOR2_X1 U2849 ( .A(n499), .B(n366), .ZN(n2683) );
  XNOR2_X1 U2850 ( .A(n499), .B(n3574), .ZN(n2749) );
  XNOR2_X1 U2851 ( .A(n499), .B(n324), .ZN(n3145) );
  XNOR2_X1 U2852 ( .A(n499), .B(n330), .ZN(n3079) );
  XNOR2_X1 U2853 ( .A(n499), .B(n321), .ZN(n3178) );
  XNOR2_X1 U2854 ( .A(n499), .B(n345), .ZN(n2914) );
  XNOR2_X1 U2855 ( .A(n499), .B(n363), .ZN(n2716) );
  XNOR2_X1 U2856 ( .A(n499), .B(n354), .ZN(n2815) );
  XNOR2_X1 U2857 ( .A(n499), .B(n327), .ZN(n3112) );
  XNOR2_X1 U2858 ( .A(n499), .B(n348), .ZN(n2881) );
  XNOR2_X1 U2859 ( .A(n499), .B(n339), .ZN(n2980) );
  XNOR2_X1 U2860 ( .A(n499), .B(n351), .ZN(n2848) );
  XNOR2_X1 U2861 ( .A(n499), .B(n342), .ZN(n2947) );
  INV_X1 U2862 ( .A(n501), .ZN(n2651) );
  XNOR2_X1 U2863 ( .A(n501), .B(n327), .ZN(n3111) );
  XNOR2_X1 U2864 ( .A(n501), .B(n357), .ZN(n2781) );
  XNOR2_X1 U2865 ( .A(n501), .B(n366), .ZN(n2682) );
  XNOR2_X1 U2866 ( .A(n501), .B(n324), .ZN(n3144) );
  XNOR2_X1 U2867 ( .A(n501), .B(n321), .ZN(n3177) );
  XNOR2_X1 U2868 ( .A(n501), .B(n330), .ZN(n3078) );
  XNOR2_X1 U2869 ( .A(n501), .B(n351), .ZN(n2847) );
  XNOR2_X1 U2870 ( .A(n501), .B(n345), .ZN(n2913) );
  XNOR2_X1 U2871 ( .A(n501), .B(n363), .ZN(n2715) );
  XNOR2_X1 U2872 ( .A(n501), .B(n3574), .ZN(n2748) );
  XNOR2_X1 U2873 ( .A(n501), .B(n354), .ZN(n2814) );
  XNOR2_X1 U2874 ( .A(n501), .B(n348), .ZN(n2880) );
  XNOR2_X1 U2875 ( .A(n501), .B(n339), .ZN(n2979) );
  XNOR2_X1 U2876 ( .A(n501), .B(n3554), .ZN(n3045) );
  XNOR2_X1 U2877 ( .A(n501), .B(n342), .ZN(n2946) );
  INV_X1 U2878 ( .A(n497), .ZN(n2653) );
  XNOR2_X1 U2879 ( .A(n497), .B(n3574), .ZN(n2750) );
  XNOR2_X1 U2880 ( .A(n497), .B(n324), .ZN(n3146) );
  XNOR2_X1 U2881 ( .A(n497), .B(n330), .ZN(n3080) );
  XNOR2_X1 U2882 ( .A(n497), .B(n321), .ZN(n3179) );
  XNOR2_X1 U2883 ( .A(n497), .B(n366), .ZN(n2684) );
  XNOR2_X1 U2884 ( .A(n497), .B(n357), .ZN(n2783) );
  XNOR2_X1 U2885 ( .A(n497), .B(n363), .ZN(n2717) );
  XNOR2_X1 U2886 ( .A(n497), .B(n348), .ZN(n2882) );
  XNOR2_X1 U2887 ( .A(n497), .B(n327), .ZN(n3113) );
  XNOR2_X1 U2888 ( .A(n497), .B(n339), .ZN(n2981) );
  XNOR2_X1 U2889 ( .A(n497), .B(n342), .ZN(n2948) );
  XNOR2_X1 U2890 ( .A(n497), .B(n336), .ZN(n3014) );
  XNOR2_X1 U2891 ( .A(n497), .B(n345), .ZN(n2915) );
  XNOR2_X1 U2892 ( .A(n497), .B(n351), .ZN(n2849) );
  XNOR2_X1 U2893 ( .A(n497), .B(n354), .ZN(n2816) );
  INV_X1 U2894 ( .A(n495), .ZN(n2654) );
  XNOR2_X1 U2895 ( .A(n495), .B(n3574), .ZN(n2751) );
  XNOR2_X1 U2896 ( .A(n495), .B(n330), .ZN(n3081) );
  XNOR2_X1 U2897 ( .A(n495), .B(n363), .ZN(n2718) );
  XNOR2_X1 U2898 ( .A(n495), .B(n321), .ZN(n3180) );
  XNOR2_X1 U2899 ( .A(n495), .B(n3554), .ZN(n3048) );
  XNOR2_X1 U2900 ( .A(n495), .B(n324), .ZN(n3147) );
  XNOR2_X1 U2901 ( .A(n495), .B(n348), .ZN(n2883) );
  XNOR2_X1 U2902 ( .A(n495), .B(n351), .ZN(n2850) );
  XNOR2_X1 U2903 ( .A(n495), .B(n366), .ZN(n2685) );
  XNOR2_X1 U2904 ( .A(n495), .B(n357), .ZN(n2784) );
  XNOR2_X1 U2905 ( .A(n495), .B(n336), .ZN(n3015) );
  XNOR2_X1 U2906 ( .A(n495), .B(n345), .ZN(n2916) );
  XNOR2_X1 U2907 ( .A(n495), .B(n339), .ZN(n2982) );
  XNOR2_X1 U2908 ( .A(n495), .B(n327), .ZN(n3114) );
  XNOR2_X1 U2909 ( .A(n495), .B(n342), .ZN(n2949) );
  XNOR2_X1 U2910 ( .A(n495), .B(n354), .ZN(n2817) );
  XNOR2_X1 U2911 ( .A(n491), .B(n3559), .ZN(n3050) );
  INV_X1 U2912 ( .A(n491), .ZN(n2656) );
  XNOR2_X1 U2913 ( .A(n491), .B(n321), .ZN(n3182) );
  XNOR2_X1 U2914 ( .A(n491), .B(n363), .ZN(n2720) );
  XNOR2_X1 U2915 ( .A(n491), .B(n351), .ZN(n2852) );
  XNOR2_X1 U2916 ( .A(n491), .B(n327), .ZN(n3116) );
  XNOR2_X1 U2917 ( .A(n491), .B(n336), .ZN(n3017) );
  XNOR2_X1 U2918 ( .A(n491), .B(n330), .ZN(n3083) );
  XNOR2_X1 U2919 ( .A(n491), .B(n366), .ZN(n2687) );
  XNOR2_X1 U2920 ( .A(n491), .B(n342), .ZN(n2951) );
  XNOR2_X1 U2921 ( .A(n491), .B(n324), .ZN(n3149) );
  XNOR2_X1 U2922 ( .A(n491), .B(n348), .ZN(n2885) );
  XNOR2_X1 U2923 ( .A(n491), .B(n345), .ZN(n2918) );
  XNOR2_X1 U2924 ( .A(n491), .B(n357), .ZN(n2786) );
  XNOR2_X1 U2925 ( .A(n491), .B(n354), .ZN(n2819) );
  XNOR2_X1 U2926 ( .A(n491), .B(n360), .ZN(n2753) );
  XNOR2_X1 U2927 ( .A(n491), .B(n339), .ZN(n2984) );
  INV_X1 U2928 ( .A(n493), .ZN(n2655) );
  XNOR2_X1 U2929 ( .A(n493), .B(n321), .ZN(n3181) );
  XNOR2_X1 U2930 ( .A(n493), .B(n363), .ZN(n2719) );
  XNOR2_X1 U2931 ( .A(n493), .B(n3574), .ZN(n2752) );
  XNOR2_X1 U2932 ( .A(n493), .B(n336), .ZN(n3016) );
  XNOR2_X1 U2933 ( .A(n493), .B(n351), .ZN(n2851) );
  XNOR2_X1 U2934 ( .A(n493), .B(n324), .ZN(n3148) );
  XNOR2_X1 U2935 ( .A(n493), .B(n3554), .ZN(n3049) );
  XNOR2_X1 U2936 ( .A(n493), .B(n330), .ZN(n3082) );
  XNOR2_X1 U2937 ( .A(n493), .B(n366), .ZN(n2686) );
  XNOR2_X1 U2938 ( .A(n493), .B(n357), .ZN(n2785) );
  XNOR2_X1 U2939 ( .A(n493), .B(n327), .ZN(n3115) );
  XNOR2_X1 U2940 ( .A(n493), .B(n348), .ZN(n2884) );
  XNOR2_X1 U2941 ( .A(n493), .B(n339), .ZN(n2983) );
  XNOR2_X1 U2942 ( .A(n493), .B(n342), .ZN(n2950) );
  XNOR2_X1 U2943 ( .A(n493), .B(n345), .ZN(n2917) );
  XNOR2_X1 U2944 ( .A(n493), .B(n354), .ZN(n2818) );
  INV_X1 U2945 ( .A(n489), .ZN(n2657) );
  XNOR2_X1 U2946 ( .A(n489), .B(n3554), .ZN(n3051) );
  XNOR2_X1 U2947 ( .A(n489), .B(n366), .ZN(n2688) );
  XNOR2_X1 U2948 ( .A(n489), .B(n330), .ZN(n3084) );
  XNOR2_X1 U2949 ( .A(n489), .B(n321), .ZN(n3183) );
  XNOR2_X1 U2950 ( .A(n489), .B(n324), .ZN(n3150) );
  XNOR2_X1 U2951 ( .A(n489), .B(n327), .ZN(n3117) );
  XNOR2_X1 U2952 ( .A(n489), .B(n363), .ZN(n2721) );
  XNOR2_X1 U2953 ( .A(n489), .B(n354), .ZN(n2820) );
  XNOR2_X1 U2954 ( .A(n489), .B(n3574), .ZN(n2754) );
  XNOR2_X1 U2955 ( .A(n489), .B(n348), .ZN(n2886) );
  XNOR2_X1 U2956 ( .A(n489), .B(n342), .ZN(n2952) );
  XNOR2_X1 U2957 ( .A(n489), .B(n345), .ZN(n2919) );
  XNOR2_X1 U2958 ( .A(n489), .B(n339), .ZN(n2985) );
  XNOR2_X1 U2959 ( .A(n489), .B(n351), .ZN(n2853) );
  INV_X1 U2960 ( .A(n487), .ZN(n2658) );
  XNOR2_X1 U2961 ( .A(n487), .B(n324), .ZN(n3151) );
  XNOR2_X1 U2962 ( .A(n487), .B(n366), .ZN(n2689) );
  XNOR2_X1 U2963 ( .A(n487), .B(n321), .ZN(n3184) );
  XNOR2_X1 U2964 ( .A(n487), .B(n330), .ZN(n3085) );
  XNOR2_X1 U2965 ( .A(n487), .B(n327), .ZN(n3118) );
  XNOR2_X1 U2966 ( .A(n487), .B(n354), .ZN(n2821) );
  XNOR2_X1 U2967 ( .A(n487), .B(n348), .ZN(n2887) );
  XNOR2_X1 U2968 ( .A(n487), .B(n363), .ZN(n2722) );
  XNOR2_X1 U2969 ( .A(n487), .B(n339), .ZN(n2986) );
  XNOR2_X1 U2970 ( .A(n487), .B(n345), .ZN(n2920) );
  XNOR2_X1 U2971 ( .A(n487), .B(n336), .ZN(n3019) );
  XNOR2_X1 U2972 ( .A(n487), .B(n3554), .ZN(n3052) );
  XNOR2_X1 U2973 ( .A(n487), .B(n357), .ZN(n2788) );
  XNOR2_X1 U2974 ( .A(n487), .B(n3574), .ZN(n2755) );
  XNOR2_X1 U2975 ( .A(n487), .B(n351), .ZN(n2854) );
  XNOR2_X1 U2976 ( .A(n487), .B(n342), .ZN(n2953) );
  INV_X1 U2977 ( .A(n483), .ZN(n2660) );
  XNOR2_X1 U2978 ( .A(n483), .B(n327), .ZN(n3120) );
  XNOR2_X1 U2979 ( .A(n483), .B(n3554), .ZN(n3054) );
  XNOR2_X1 U2980 ( .A(n483), .B(n321), .ZN(n3186) );
  XNOR2_X1 U2981 ( .A(n483), .B(n363), .ZN(n2724) );
  XNOR2_X1 U2982 ( .A(n483), .B(n357), .ZN(n2790) );
  XNOR2_X1 U2983 ( .A(n483), .B(n324), .ZN(n3153) );
  XNOR2_X1 U2984 ( .A(n483), .B(n366), .ZN(n2691) );
  XNOR2_X1 U2985 ( .A(n483), .B(n348), .ZN(n2889) );
  XNOR2_X1 U2986 ( .A(n483), .B(n342), .ZN(n2955) );
  XNOR2_X1 U2987 ( .A(n483), .B(n354), .ZN(n2823) );
  XNOR2_X1 U2988 ( .A(n483), .B(n339), .ZN(n2988) );
  XNOR2_X1 U2989 ( .A(n483), .B(n330), .ZN(n3087) );
  XNOR2_X1 U2990 ( .A(n483), .B(n351), .ZN(n2856) );
  XNOR2_X1 U2991 ( .A(n483), .B(n345), .ZN(n2922) );
  XNOR2_X1 U2992 ( .A(n483), .B(n360), .ZN(n2757) );
  INV_X1 U2993 ( .A(n485), .ZN(n2659) );
  XNOR2_X1 U2994 ( .A(n485), .B(n327), .ZN(n3119) );
  XNOR2_X1 U2995 ( .A(n485), .B(n321), .ZN(n3185) );
  XNOR2_X1 U2996 ( .A(n485), .B(n363), .ZN(n2723) );
  XNOR2_X1 U2997 ( .A(n485), .B(n339), .ZN(n2987) );
  XNOR2_X1 U2998 ( .A(n485), .B(n354), .ZN(n2822) );
  XNOR2_X1 U2999 ( .A(n485), .B(n324), .ZN(n3152) );
  XNOR2_X1 U3000 ( .A(n485), .B(n366), .ZN(n2690) );
  XNOR2_X1 U3001 ( .A(n485), .B(n348), .ZN(n2888) );
  XNOR2_X1 U3002 ( .A(n485), .B(n3554), .ZN(n3053) );
  XNOR2_X1 U3003 ( .A(n485), .B(n357), .ZN(n2789) );
  XNOR2_X1 U3004 ( .A(n485), .B(n3574), .ZN(n2756) );
  XNOR2_X1 U3005 ( .A(n485), .B(n330), .ZN(n3086) );
  XNOR2_X1 U3006 ( .A(n485), .B(n351), .ZN(n2855) );
  XNOR2_X1 U3007 ( .A(n485), .B(n345), .ZN(n2921) );
  XNOR2_X1 U3008 ( .A(n485), .B(n342), .ZN(n2954) );
  INV_X1 U3009 ( .A(n481), .ZN(n2661) );
  XNOR2_X1 U3010 ( .A(n481), .B(n321), .ZN(n3187) );
  XNOR2_X1 U3011 ( .A(n481), .B(n3554), .ZN(n3055) );
  XNOR2_X1 U3012 ( .A(n481), .B(n324), .ZN(n3154) );
  XNOR2_X1 U3013 ( .A(n481), .B(n330), .ZN(n3088) );
  XNOR2_X1 U3014 ( .A(n481), .B(n363), .ZN(n2725) );
  XNOR2_X1 U3015 ( .A(n481), .B(n351), .ZN(n2857) );
  XNOR2_X1 U3016 ( .A(n481), .B(n366), .ZN(n2692) );
  XNOR2_X1 U3017 ( .A(n481), .B(n327), .ZN(n3121) );
  XNOR2_X1 U3018 ( .A(n481), .B(n357), .ZN(n2791) );
  XNOR2_X1 U3019 ( .A(n481), .B(n342), .ZN(n2956) );
  XNOR2_X1 U3020 ( .A(n481), .B(n345), .ZN(n2923) );
  XNOR2_X1 U3021 ( .A(n481), .B(n336), .ZN(n3022) );
  XNOR2_X1 U3022 ( .A(n481), .B(n360), .ZN(n2758) );
  XNOR2_X1 U3023 ( .A(n481), .B(n354), .ZN(n2824) );
  XNOR2_X1 U3024 ( .A(n481), .B(n339), .ZN(n2989) );
  XNOR2_X1 U3025 ( .A(n481), .B(n348), .ZN(n2890) );
  INV_X1 U3026 ( .A(n479), .ZN(n2662) );
  XNOR2_X1 U3027 ( .A(n479), .B(n321), .ZN(n3188) );
  XNOR2_X1 U3028 ( .A(n479), .B(n324), .ZN(n3155) );
  XNOR2_X1 U3029 ( .A(n479), .B(n345), .ZN(n2924) );
  XNOR2_X1 U3030 ( .A(n479), .B(n327), .ZN(n3122) );
  XNOR2_X1 U3031 ( .A(n479), .B(n330), .ZN(n3089) );
  XNOR2_X1 U3032 ( .A(n479), .B(n336), .ZN(n3023) );
  XNOR2_X1 U3033 ( .A(n479), .B(n339), .ZN(n2990) );
  XNOR2_X1 U3034 ( .A(n479), .B(n342), .ZN(n2957) );
  XNOR2_X1 U3035 ( .A(n479), .B(n351), .ZN(n2858) );
  XNOR2_X1 U3036 ( .A(n479), .B(n354), .ZN(n2825) );
  XNOR2_X1 U3037 ( .A(n479), .B(n3554), .ZN(n3056) );
  XNOR2_X1 U3038 ( .A(n479), .B(n360), .ZN(n2759) );
  XNOR2_X1 U3039 ( .A(n479), .B(n357), .ZN(n2792) );
  XNOR2_X1 U3040 ( .A(n479), .B(n348), .ZN(n2891) );
  XNOR2_X1 U3041 ( .A(n479), .B(n363), .ZN(n2726) );
  XNOR2_X1 U3042 ( .A(n479), .B(n366), .ZN(n2693) );
  XNOR2_X1 U3043 ( .A(n475), .B(n321), .ZN(n3190) );
  INV_X1 U3044 ( .A(n475), .ZN(n2664) );
  XNOR2_X1 U3045 ( .A(n475), .B(n324), .ZN(n3157) );
  XNOR2_X1 U3046 ( .A(n475), .B(n327), .ZN(n3124) );
  XNOR2_X1 U3047 ( .A(n475), .B(n3559), .ZN(n3058) );
  XNOR2_X1 U3048 ( .A(n475), .B(n354), .ZN(n2827) );
  XNOR2_X1 U3049 ( .A(n475), .B(n339), .ZN(n2992) );
  XNOR2_X1 U3050 ( .A(n475), .B(n330), .ZN(n3091) );
  XNOR2_X1 U3051 ( .A(n475), .B(n342), .ZN(n2959) );
  XNOR2_X1 U3052 ( .A(n475), .B(n345), .ZN(n2926) );
  XNOR2_X1 U3053 ( .A(n475), .B(n348), .ZN(n2893) );
  XNOR2_X1 U3054 ( .A(n475), .B(n357), .ZN(n2794) );
  XNOR2_X1 U3055 ( .A(n475), .B(n336), .ZN(n3025) );
  XNOR2_X1 U3056 ( .A(n475), .B(n363), .ZN(n2728) );
  XNOR2_X1 U3057 ( .A(n475), .B(n3574), .ZN(n2761) );
  XNOR2_X1 U3058 ( .A(n475), .B(n366), .ZN(n2695) );
  XNOR2_X1 U3059 ( .A(n475), .B(n351), .ZN(n2860) );
  INV_X1 U3060 ( .A(n477), .ZN(n2663) );
  XNOR2_X1 U3061 ( .A(n477), .B(n321), .ZN(n3189) );
  XNOR2_X1 U3062 ( .A(n477), .B(n324), .ZN(n3156) );
  XNOR2_X1 U3063 ( .A(n477), .B(n330), .ZN(n3090) );
  XNOR2_X1 U3064 ( .A(n477), .B(n327), .ZN(n3123) );
  XNOR2_X1 U3065 ( .A(n477), .B(n339), .ZN(n2991) );
  XNOR2_X1 U3066 ( .A(n477), .B(n354), .ZN(n2826) );
  XNOR2_X1 U3067 ( .A(n477), .B(n342), .ZN(n2958) );
  XNOR2_X1 U3068 ( .A(n477), .B(n336), .ZN(n3024) );
  XNOR2_X1 U3069 ( .A(n477), .B(n345), .ZN(n2925) );
  XNOR2_X1 U3070 ( .A(n477), .B(n3554), .ZN(n3057) );
  XNOR2_X1 U3071 ( .A(n477), .B(n348), .ZN(n2892) );
  XNOR2_X1 U3072 ( .A(n477), .B(n360), .ZN(n2760) );
  XNOR2_X1 U3073 ( .A(n477), .B(n363), .ZN(n2727) );
  XNOR2_X1 U3074 ( .A(n477), .B(n357), .ZN(n2793) );
  XNOR2_X1 U3075 ( .A(n477), .B(n366), .ZN(n2694) );
  XNOR2_X1 U3076 ( .A(n477), .B(n351), .ZN(n2859) );
  XNOR2_X1 U3077 ( .A(n473), .B(n324), .ZN(n3158) );
  INV_X1 U3078 ( .A(n473), .ZN(n2665) );
  XNOR2_X1 U3079 ( .A(n473), .B(n321), .ZN(n3191) );
  XNOR2_X1 U3080 ( .A(n473), .B(n327), .ZN(n3125) );
  XNOR2_X1 U3081 ( .A(n473), .B(n3559), .ZN(n3059) );
  XNOR2_X1 U3082 ( .A(n473), .B(n348), .ZN(n2894) );
  XNOR2_X1 U3083 ( .A(n473), .B(n345), .ZN(n2927) );
  XNOR2_X1 U3084 ( .A(n473), .B(n330), .ZN(n3092) );
  XNOR2_X1 U3085 ( .A(n473), .B(n342), .ZN(n2960) );
  XNOR2_X1 U3086 ( .A(n473), .B(n336), .ZN(n3026) );
  XNOR2_X1 U3087 ( .A(n473), .B(n357), .ZN(n2795) );
  XNOR2_X1 U3088 ( .A(n473), .B(n351), .ZN(n2861) );
  XNOR2_X1 U3089 ( .A(n473), .B(n363), .ZN(n2729) );
  XNOR2_X1 U3090 ( .A(n473), .B(n339), .ZN(n2993) );
  XNOR2_X1 U3091 ( .A(n473), .B(n3574), .ZN(n2762) );
  XNOR2_X1 U3092 ( .A(n473), .B(n366), .ZN(n2696) );
  XNOR2_X1 U3093 ( .A(n473), .B(n354), .ZN(n2828) );
  XNOR2_X1 U3094 ( .A(n471), .B(n324), .ZN(n3159) );
  INV_X1 U3095 ( .A(n471), .ZN(n2666) );
  XNOR2_X1 U3096 ( .A(n471), .B(n321), .ZN(n3192) );
  XNOR2_X1 U3097 ( .A(n471), .B(n3559), .ZN(n3060) );
  XNOR2_X1 U3098 ( .A(n471), .B(n327), .ZN(n3126) );
  XNOR2_X1 U3099 ( .A(n471), .B(n336), .ZN(n3027) );
  XNOR2_X1 U3100 ( .A(n471), .B(n330), .ZN(n3093) );
  XNOR2_X1 U3101 ( .A(n471), .B(n357), .ZN(n2796) );
  XNOR2_X1 U3102 ( .A(n471), .B(n345), .ZN(n2928) );
  XNOR2_X1 U3103 ( .A(n471), .B(n342), .ZN(n2961) );
  XNOR2_X1 U3104 ( .A(n471), .B(n360), .ZN(n2763) );
  XNOR2_X1 U3105 ( .A(n471), .B(n366), .ZN(n2697) );
  XNOR2_X1 U3106 ( .A(n471), .B(n339), .ZN(n2994) );
  XNOR2_X1 U3107 ( .A(n471), .B(n351), .ZN(n2862) );
  XNOR2_X1 U3108 ( .A(n471), .B(n348), .ZN(n2895) );
  XNOR2_X1 U3109 ( .A(n471), .B(n354), .ZN(n2829) );
  XNOR2_X1 U3110 ( .A(n471), .B(n363), .ZN(n2730) );
  XNOR2_X1 U3111 ( .A(n469), .B(n321), .ZN(n3193) );
  XNOR2_X1 U3112 ( .A(n469), .B(n3559), .ZN(n3061) );
  INV_X1 U3113 ( .A(n469), .ZN(n2667) );
  XNOR2_X1 U3114 ( .A(n469), .B(n327), .ZN(n3127) );
  XNOR2_X1 U3115 ( .A(n469), .B(n324), .ZN(n3160) );
  XNOR2_X1 U3116 ( .A(n469), .B(n3669), .ZN(n3028) );
  XNOR2_X1 U3117 ( .A(n469), .B(n360), .ZN(n2764) );
  XNOR2_X1 U3118 ( .A(n469), .B(n345), .ZN(n2929) );
  XNOR2_X1 U3119 ( .A(n469), .B(n342), .ZN(n2962) );
  XNOR2_X1 U3120 ( .A(n469), .B(n366), .ZN(n2698) );
  XNOR2_X1 U3121 ( .A(n469), .B(n339), .ZN(n2995) );
  XNOR2_X1 U3122 ( .A(n469), .B(n330), .ZN(n3094) );
  XNOR2_X1 U3123 ( .A(n469), .B(n357), .ZN(n2797) );
  XNOR2_X1 U3124 ( .A(n469), .B(n354), .ZN(n2830) );
  XNOR2_X1 U3125 ( .A(n469), .B(n348), .ZN(n2896) );
  XNOR2_X1 U3126 ( .A(n469), .B(n351), .ZN(n2863) );
  XNOR2_X1 U3127 ( .A(n469), .B(n363), .ZN(n2731) );
  XNOR2_X1 U3128 ( .A(n465), .B(n327), .ZN(n3128) );
  XNOR2_X1 U3129 ( .A(n465), .B(n321), .ZN(n3194) );
  AND2_X1 U3130 ( .A1(n465), .A2(n366), .ZN(n2093) );
  XNOR2_X1 U3131 ( .A(n465), .B(n3559), .ZN(n3062) );
  XNOR2_X1 U3132 ( .A(n465), .B(n345), .ZN(n2930) );
  XNOR2_X1 U3133 ( .A(n465), .B(n3669), .ZN(n3029) );
  XNOR2_X1 U3134 ( .A(n465), .B(n324), .ZN(n3161) );
  XNOR2_X1 U3135 ( .A(n465), .B(n3574), .ZN(n2765) );
  XNOR2_X1 U3136 ( .A(n465), .B(n342), .ZN(n2963) );
  XNOR2_X1 U3137 ( .A(n465), .B(n348), .ZN(n2897) );
  XNOR2_X1 U3138 ( .A(n465), .B(n351), .ZN(n2864) );
  XNOR2_X1 U3139 ( .A(n465), .B(n3647), .ZN(n2996) );
  XNOR2_X1 U3140 ( .A(n465), .B(n363), .ZN(n2732) );
  XNOR2_X1 U3141 ( .A(n465), .B(n330), .ZN(n3095) );
  XNOR2_X1 U3142 ( .A(n465), .B(n354), .ZN(n2831) );
  XNOR2_X1 U3143 ( .A(n465), .B(n366), .ZN(n2699) );
  XNOR2_X1 U3144 ( .A(n465), .B(n357), .ZN(n2798) );
  INV_X2 U3145 ( .A(n363), .ZN(n3512) );
  INV_X1 U3146 ( .A(n824), .ZN(n822) );
  XNOR2_X2 U3147 ( .A(n3737), .B(n330), .ZN(n3577) );
  NAND2_X1 U3148 ( .A1(n1670), .A2(n1697), .ZN(n820) );
  NOR2_X1 U3149 ( .A1(n819), .A2(n824), .ZN(n817) );
  NOR2_X1 U3150 ( .A1(n1377), .A2(n1402), .ZN(n3409) );
  NOR2_X1 U3151 ( .A1(n1377), .A2(n1402), .ZN(n769) );
  INV_X1 U3152 ( .A(n3554), .ZN(n3558) );
  NAND2_X1 U3153 ( .A1(a[22]), .A2(n3615), .ZN(n3616) );
  INV_X2 U3154 ( .A(n351), .ZN(n3615) );
  OAI21_X2 U3155 ( .B1(n819), .B2(n825), .A(n820), .ZN(n818) );
  OAI22_X1 U3156 ( .A1(n3475), .A2(n2860), .B1(n2859), .B2(n3672), .ZN(n2292)
         );
  XNOR2_X1 U3157 ( .A(n3415), .B(n348), .ZN(n3234) );
  XOR2_X2 U3158 ( .A(n1645), .B(n3411), .Z(n1614) );
  BUF_X1 U3159 ( .A(n814), .Z(n3410) );
  INV_X2 U3160 ( .A(n333), .ZN(n3553) );
  AND2_X2 U3161 ( .A1(n3229), .A2(n3521), .ZN(n3742) );
  INV_X1 U3162 ( .A(n907), .ZN(n1026) );
  OAI21_X2 U3163 ( .B1(n907), .B2(n913), .A(n908), .ZN(n906) );
  XOR2_X1 U3164 ( .A(n1618), .B(n1620), .Z(n3411) );
  NAND2_X1 U3165 ( .A1(n1645), .A2(n1618), .ZN(n3412) );
  NAND2_X1 U3166 ( .A1(n1645), .A2(n1620), .ZN(n3413) );
  NAND2_X1 U3167 ( .A1(n1618), .A2(n1620), .ZN(n3414) );
  NAND3_X1 U3168 ( .A1(n3412), .A2(n3414), .A3(n3413), .ZN(n1613) );
  NAND2_X1 U3169 ( .A1(a[18]), .A2(n345), .ZN(n3417) );
  NAND2_X1 U3170 ( .A1(n3415), .A2(n3416), .ZN(n3418) );
  NAND2_X1 U3171 ( .A1(n3417), .A2(n3418), .ZN(n3550) );
  INV_X1 U3172 ( .A(a[18]), .ZN(n3415) );
  INV_X1 U3173 ( .A(n345), .ZN(n3416) );
  INV_X1 U3174 ( .A(n3550), .ZN(n3696) );
  XNOR2_X1 U3175 ( .A(n3745), .B(n366), .ZN(n3228) );
  INV_X1 U3176 ( .A(n847), .ZN(n845) );
  OAI21_X2 U3177 ( .B1(n877), .B2(n857), .A(n858), .ZN(n856) );
  OAI22_X1 U3178 ( .A1(n3693), .A2(n3012), .B1(n3011), .B2(n3566), .ZN(n2449)
         );
  BUF_X1 U3179 ( .A(n3628), .Z(n3419) );
  NAND2_X1 U3180 ( .A1(a[2]), .A2(n3421), .ZN(n3422) );
  NAND2_X1 U3181 ( .A1(n3420), .A2(n324), .ZN(n3423) );
  NAND2_X1 U3182 ( .A1(n3422), .A2(n3423), .ZN(n3242) );
  INV_X1 U3183 ( .A(a[2]), .ZN(n3420) );
  INV_X1 U3184 ( .A(n324), .ZN(n3421) );
  AND2_X1 U3185 ( .A1(n3242), .A2(n3648), .ZN(n3750) );
  NOR2_X1 U3186 ( .A1(n727), .A2(n613), .ZN(n611) );
  INV_X1 U3187 ( .A(n727), .ZN(n725) );
  NAND2_X1 U3188 ( .A1(n752), .A2(n729), .ZN(n727) );
  NAND2_X1 U3189 ( .A1(n1259), .A2(n1280), .ZN(n736) );
  XNOR2_X1 U3190 ( .A(n3737), .B(n3290), .ZN(n3424) );
  INV_X4 U3191 ( .A(n327), .ZN(n3290) );
  OAI21_X2 U3192 ( .B1(n3556), .B2(n804), .A(n801), .ZN(n799) );
  NAND2_X2 U3193 ( .A1(n3605), .A2(n3606), .ZN(n3706) );
  XNOR2_X1 U3194 ( .A(n3614), .B(n354), .ZN(n3232) );
  XOR2_X1 U3195 ( .A(n2279), .B(n2119), .Z(n3425) );
  XOR2_X1 U3196 ( .A(n2439), .B(n3425), .Z(n1425) );
  NAND2_X1 U3197 ( .A1(n2439), .A2(n2279), .ZN(n3426) );
  NAND2_X1 U3198 ( .A1(n2439), .A2(n2119), .ZN(n3427) );
  NAND2_X1 U3199 ( .A1(n2279), .A2(n2119), .ZN(n3428) );
  NAND3_X1 U3200 ( .A1(n3426), .A2(n3428), .A3(n3427), .ZN(n1424) );
  AOI21_X1 U3201 ( .B1(n753), .B2(n729), .A(n730), .ZN(n3429) );
  OR2_X1 U3202 ( .A1(n3551), .A2(n3002), .ZN(n3430) );
  OR2_X1 U3203 ( .A1(n3001), .A2(n3566), .ZN(n3431) );
  NAND2_X1 U3204 ( .A1(n3430), .A2(n3431), .ZN(n2439) );
  OAI22_X1 U3205 ( .A1(n3475), .A2(n2847), .B1(n2846), .B2(n3673), .ZN(n2279)
         );
  AOI21_X1 U3206 ( .B1(n753), .B2(n729), .A(n730), .ZN(n728) );
  XNOR2_X1 U3207 ( .A(n521), .B(n336), .ZN(n3002) );
  XNOR2_X1 U3208 ( .A(n523), .B(n336), .ZN(n3001) );
  XNOR2_X1 U3209 ( .A(n3749), .B(n327), .ZN(n3241) );
  INV_X1 U3210 ( .A(n3664), .ZN(n3432) );
  XNOR2_X1 U3211 ( .A(n1726), .B(n3433), .ZN(n1724) );
  XNOR2_X1 U3212 ( .A(n1751), .B(n1728), .ZN(n3433) );
  XOR2_X1 U3213 ( .A(n2458), .B(n2586), .Z(n3434) );
  XOR2_X1 U3214 ( .A(n3434), .B(n2554), .Z(n1910) );
  XOR2_X1 U3215 ( .A(n1927), .B(n1912), .Z(n3435) );
  XOR2_X1 U3216 ( .A(n3435), .B(n1910), .Z(n1906) );
  NAND2_X1 U3217 ( .A1(n2458), .A2(n2586), .ZN(n3436) );
  NAND2_X1 U3218 ( .A1(n2458), .A2(n2554), .ZN(n3437) );
  NAND2_X1 U3219 ( .A1(n2586), .A2(n2554), .ZN(n3438) );
  NAND3_X1 U3220 ( .A1(n3436), .A2(n3437), .A3(n3438), .ZN(n1909) );
  NAND2_X1 U3221 ( .A1(n1927), .A2(n1912), .ZN(n3439) );
  NAND2_X1 U3222 ( .A1(n1927), .A2(n1910), .ZN(n3440) );
  NAND2_X1 U3223 ( .A1(n1912), .A2(n1910), .ZN(n3441) );
  NAND3_X1 U3224 ( .A1(n3439), .A2(n3440), .A3(n3441), .ZN(n1905) );
  BUF_X1 U3225 ( .A(n856), .Z(n3442) );
  OR2_X1 U3226 ( .A1(n3552), .A2(n3021), .ZN(n3443) );
  OR2_X1 U3227 ( .A1(n3020), .A2(n3567), .ZN(n3444) );
  NAND2_X1 U3228 ( .A1(n3443), .A2(n3444), .ZN(n2458) );
  XNOR2_X1 U3229 ( .A(n483), .B(n336), .ZN(n3021) );
  XNOR2_X1 U3230 ( .A(n485), .B(n336), .ZN(n3020) );
  FA_X1 U3231 ( .A(n1643), .B(n1616), .CI(n1614), .S(n3445) );
  INV_X1 U3232 ( .A(n696), .ZN(n992) );
  OAI21_X1 U3233 ( .B1(n696), .B2(n700), .A(n697), .ZN(n695) );
  NAND2_X1 U3234 ( .A1(n1167), .A2(n1182), .ZN(n697) );
  OAI22_X1 U3235 ( .A1(n452), .A2(n2817), .B1(n2816), .B2(n402), .ZN(n2248) );
  INV_X4 U3236 ( .A(n3680), .ZN(n437) );
  NAND2_X2 U3237 ( .A1(n3739), .A2(n336), .ZN(n3621) );
  INV_X4 U3238 ( .A(a[12]), .ZN(n3739) );
  NOR2_X1 U3239 ( .A1(n883), .A2(n880), .ZN(n878) );
  OAI22_X1 U3240 ( .A1(n428), .A2(n3087), .B1(n3086), .B2(n3664), .ZN(n2526)
         );
  OAI21_X1 U3241 ( .B1(n884), .B2(n880), .A(n881), .ZN(n879) );
  AND2_X2 U3242 ( .A1(n3241), .A2(n3532), .ZN(n3684) );
  INV_X1 U3243 ( .A(n758), .ZN(n3446) );
  OR2_X1 U3244 ( .A1(n1327), .A2(n1350), .ZN(n3447) );
  OAI22_X1 U3245 ( .A1(n419), .A2(n3189), .B1(n3188), .B2(n3511), .ZN(n2631)
         );
  OAI22_X1 U3246 ( .A1(n419), .A2(n3188), .B1(n3187), .B2(n3511), .ZN(n2630)
         );
  OAI22_X1 U3247 ( .A1(n419), .A2(n3178), .B1(n3177), .B2(n3511), .ZN(n2620)
         );
  OAI22_X1 U3248 ( .A1(n419), .A2(n3187), .B1(n3186), .B2(n3511), .ZN(n2629)
         );
  OAI22_X1 U3249 ( .A1(n419), .A2(n3185), .B1(n3184), .B2(n3511), .ZN(n2627)
         );
  OAI22_X1 U3250 ( .A1(n419), .A2(n3181), .B1(n3180), .B2(n3511), .ZN(n2623)
         );
  OAI22_X1 U3251 ( .A1(n419), .A2(n3174), .B1(n3173), .B2(n3511), .ZN(n2616)
         );
  OAI22_X1 U3252 ( .A1(n419), .A2(n3183), .B1(n3182), .B2(n3511), .ZN(n2625)
         );
  OAI22_X1 U3253 ( .A1(n419), .A2(n3182), .B1(n3181), .B2(n3511), .ZN(n2624)
         );
  OAI22_X1 U3254 ( .A1(n419), .A2(n3163), .B1(n3292), .B2(n3511), .ZN(n2605)
         );
  OAI22_X1 U3255 ( .A1(n419), .A2(n3184), .B1(n3183), .B2(n3511), .ZN(n2626)
         );
  OAI22_X1 U3256 ( .A1(n419), .A2(n3169), .B1(n3168), .B2(n3511), .ZN(n2611)
         );
  OAI22_X1 U3257 ( .A1(n419), .A2(n3179), .B1(n3178), .B2(n3511), .ZN(n2621)
         );
  OAI22_X1 U3258 ( .A1(n419), .A2(n3172), .B1(n3171), .B2(n3511), .ZN(n2614)
         );
  OAI22_X1 U3259 ( .A1(n419), .A2(n3176), .B1(n3175), .B2(n3511), .ZN(n2618)
         );
  OAI22_X1 U3260 ( .A1(n419), .A2(n3173), .B1(n3172), .B2(n3511), .ZN(n2615)
         );
  OAI22_X1 U3261 ( .A1(n419), .A2(n3177), .B1(n3176), .B2(n3511), .ZN(n2619)
         );
  OAI22_X1 U3262 ( .A1(n419), .A2(n3168), .B1(n3167), .B2(n3511), .ZN(n2610)
         );
  OAI22_X1 U3263 ( .A1(n419), .A2(n3180), .B1(n3179), .B2(n3511), .ZN(n2622)
         );
  OAI22_X1 U3264 ( .A1(n419), .A2(n3170), .B1(n3169), .B2(n3511), .ZN(n2612)
         );
  OAI22_X1 U3265 ( .A1(n419), .A2(n3167), .B1(n3166), .B2(n3511), .ZN(n2609)
         );
  OAI22_X1 U3266 ( .A1(n419), .A2(n3171), .B1(n3170), .B2(n3511), .ZN(n2613)
         );
  NAND2_X1 U3267 ( .A1(n1798), .A2(n1819), .ZN(n850) );
  NOR2_X1 U3268 ( .A1(n1798), .A2(n1819), .ZN(n849) );
  OAI22_X1 U3269 ( .A1(n3683), .A2(n2896), .B1(n2895), .B2(n396), .ZN(n2329)
         );
  XOR2_X1 U3270 ( .A(n2408), .B(n2248), .Z(n3448) );
  XOR2_X2 U3271 ( .A(n2440), .B(n3448), .Z(n1451) );
  XOR2_X1 U3272 ( .A(n1457), .B(n1449), .Z(n3449) );
  XOR2_X1 U3273 ( .A(n3449), .B(n1451), .Z(n1443) );
  NAND2_X1 U3274 ( .A1(n2408), .A2(n2248), .ZN(n3450) );
  NAND2_X1 U3275 ( .A1(n2408), .A2(n2440), .ZN(n3451) );
  NAND2_X4 U3276 ( .A1(n2248), .A2(n2440), .ZN(n3452) );
  NAND3_X1 U3277 ( .A1(n3450), .A2(n3451), .A3(n3452), .ZN(n1450) );
  NAND2_X1 U3278 ( .A1(n1457), .A2(n1449), .ZN(n3453) );
  NAND2_X1 U3279 ( .A1(n1457), .A2(n1451), .ZN(n3454) );
  NAND2_X1 U3280 ( .A1(n1449), .A2(n1451), .ZN(n3455) );
  NAND3_X1 U3281 ( .A1(n3453), .A2(n3454), .A3(n3455), .ZN(n1442) );
  XNOR2_X1 U3282 ( .A(n507), .B(n3554), .ZN(n3042) );
  XNOR2_X1 U3283 ( .A(n499), .B(n333), .ZN(n3046) );
  XNOR2_X1 U3284 ( .A(n497), .B(n333), .ZN(n3047) );
  XNOR2_X1 U3285 ( .A(n511), .B(n333), .ZN(n3040) );
  XNOR2_X1 U3286 ( .A(n525), .B(n333), .ZN(n3033) );
  XNOR2_X1 U3287 ( .A(n527), .B(n333), .ZN(n3032) );
  OAI22_X1 U3288 ( .A1(n437), .A2(n2975), .B1(n2974), .B2(n3571), .ZN(n2411)
         );
  OAI22_X1 U3289 ( .A1(n437), .A2(n2988), .B1(n2987), .B2(n3571), .ZN(n2424)
         );
  OAI22_X1 U3290 ( .A1(n437), .A2(n2992), .B1(n2991), .B2(n3571), .ZN(n2428)
         );
  OAI22_X1 U3291 ( .A1(n437), .A2(n2968), .B1(n2967), .B2(n3571), .ZN(n2404)
         );
  OAI22_X1 U3292 ( .A1(n437), .A2(n2977), .B1(n2976), .B2(n3571), .ZN(n2413)
         );
  OAI22_X1 U3293 ( .A1(n437), .A2(n2987), .B1(n2986), .B2(n3571), .ZN(n2423)
         );
  OAI22_X1 U3294 ( .A1(n437), .A2(n2973), .B1(n2972), .B2(n3571), .ZN(n2409)
         );
  OAI22_X1 U3295 ( .A1(n437), .A2(n2967), .B1(n2966), .B2(n3571), .ZN(n2403)
         );
  OAI22_X1 U3296 ( .A1(n437), .A2(n2981), .B1(n2980), .B2(n3571), .ZN(n2417)
         );
  OAI22_X1 U3297 ( .A1(n437), .A2(n2980), .B1(n2979), .B2(n3571), .ZN(n2416)
         );
  OAI22_X1 U3298 ( .A1(n437), .A2(n2984), .B1(n2983), .B2(n3571), .ZN(n2420)
         );
  OAI22_X1 U3299 ( .A1(n437), .A2(n2979), .B1(n2978), .B2(n3571), .ZN(n2415)
         );
  OAI22_X1 U3300 ( .A1(n437), .A2(n2965), .B1(n3571), .B2(n3286), .ZN(n2401)
         );
  OAI22_X1 U3301 ( .A1(n437), .A2(n2978), .B1(n2977), .B2(n3571), .ZN(n2414)
         );
  OAI22_X1 U3302 ( .A1(n437), .A2(n2985), .B1(n2984), .B2(n3571), .ZN(n2421)
         );
  OAI22_X1 U3303 ( .A1(n437), .A2(n2970), .B1(n2969), .B2(n3571), .ZN(n2406)
         );
  OAI22_X1 U3304 ( .A1(n437), .A2(n2972), .B1(n2971), .B2(n3571), .ZN(n2408)
         );
  AND2_X2 U3305 ( .A1(n3237), .A2(n387), .ZN(n3680) );
  BUF_X1 U3306 ( .A(n772), .Z(n3456) );
  XNOR2_X1 U3307 ( .A(n1491), .B(n3457), .ZN(n1489) );
  XNOR2_X1 U3308 ( .A(n1520), .B(n1493), .ZN(n3457) );
  BUF_X1 U3309 ( .A(n3607), .Z(n3458) );
  BUF_X8 U3310 ( .A(n3607), .Z(n3459) );
  OR2_X2 U3311 ( .A1(n3546), .A2(n3700), .ZN(n3607) );
  INV_X8 U3312 ( .A(n3736), .ZN(n446) );
  OAI22_X1 U3313 ( .A1(n3602), .A2(n3056), .B1(n3055), .B2(n381), .ZN(n2494)
         );
  OAI22_X1 U3314 ( .A1(n3602), .A2(n3051), .B1(n3050), .B2(n381), .ZN(n2489)
         );
  OAI22_X1 U3315 ( .A1(n3602), .A2(n3042), .B1(n3041), .B2(n381), .ZN(n2480)
         );
  OAI22_X1 U3316 ( .A1(n3602), .A2(n3062), .B1(n3061), .B2(n381), .ZN(n2500)
         );
  OAI22_X1 U3317 ( .A1(n3602), .A2(n3061), .B1(n3060), .B2(n381), .ZN(n2499)
         );
  OAI22_X1 U3318 ( .A1(n3602), .A2(n3054), .B1(n3053), .B2(n381), .ZN(n2492)
         );
  OAI22_X1 U3319 ( .A1(n3602), .A2(n3057), .B1(n3056), .B2(n381), .ZN(n2495)
         );
  OAI22_X1 U3320 ( .A1(n3602), .A2(n3039), .B1(n3038), .B2(n381), .ZN(n2477)
         );
  OAI22_X1 U3321 ( .A1(n3602), .A2(n3046), .B1(n3045), .B2(n381), .ZN(n2484)
         );
  OAI22_X1 U3322 ( .A1(n3602), .A2(n3033), .B1(n3032), .B2(n381), .ZN(n2471)
         );
  OR2_X2 U3323 ( .A1(n1774), .A2(n1797), .ZN(n3460) );
  OAI22_X1 U3324 ( .A1(n419), .A2(n3175), .B1(n3174), .B2(n3511), .ZN(n2617)
         );
  NOR2_X2 U3325 ( .A1(n861), .A2(n864), .ZN(n859) );
  INV_X2 U3326 ( .A(n416), .ZN(n3461) );
  INV_X8 U3327 ( .A(n3461), .ZN(n3462) );
  XOR2_X1 U3328 ( .A(n2443), .B(n2315), .Z(n3463) );
  XOR2_X1 U3329 ( .A(n3463), .B(n2347), .Z(n1539) );
  XOR2_X1 U3330 ( .A(n1547), .B(n1572), .Z(n3464) );
  XOR2_X1 U3331 ( .A(n3464), .B(n1539), .Z(n1533) );
  NAND2_X1 U3332 ( .A1(n2315), .A2(n2443), .ZN(n3465) );
  NAND2_X1 U3333 ( .A1(n2315), .A2(n2347), .ZN(n3466) );
  NAND2_X1 U3334 ( .A1(n2443), .A2(n2347), .ZN(n3467) );
  NAND3_X1 U3335 ( .A1(n3465), .A2(n3466), .A3(n3467), .ZN(n1538) );
  NAND2_X1 U3336 ( .A1(n1547), .A2(n1572), .ZN(n3468) );
  NAND2_X1 U3337 ( .A1(n1547), .A2(n1539), .ZN(n3469) );
  NAND2_X1 U3338 ( .A1(n1572), .A2(n1539), .ZN(n3470) );
  NAND3_X1 U3339 ( .A1(n3468), .A2(n3469), .A3(n3470), .ZN(n1532) );
  INV_X8 U3340 ( .A(n3662), .ZN(n3471) );
  AND2_X4 U3341 ( .A1(n3231), .A2(n3650), .ZN(n3662) );
  INV_X4 U3342 ( .A(n3662), .ZN(n455) );
  AOI21_X2 U3343 ( .B1(n997), .B2(n3509), .A(n734), .ZN(n732) );
  BUF_X1 U3344 ( .A(n773), .Z(n3473) );
  NAND2_X1 U3345 ( .A1(n1489), .A2(n1518), .ZN(n789) );
  INV_X2 U3346 ( .A(n3587), .ZN(n3475) );
  INV_X4 U3347 ( .A(n3587), .ZN(n3474) );
  INV_X1 U3348 ( .A(n399), .ZN(n3476) );
  INV_X1 U3349 ( .A(n3587), .ZN(n449) );
  INV_X2 U3350 ( .A(n3740), .ZN(n399) );
  XNOR2_X1 U3351 ( .A(n779), .B(n558), .ZN(product[37]) );
  XOR2_X1 U3352 ( .A(n782), .B(n559), .Z(product[36]) );
  NOR2_X4 U3353 ( .A1(n1862), .A2(n1881), .ZN(n869) );
  XOR2_X1 U3354 ( .A(n1699), .B(n1674), .Z(n3477) );
  XOR2_X1 U3355 ( .A(n1672), .B(n3477), .Z(n1670) );
  NAND2_X1 U3356 ( .A1(n1672), .A2(n1699), .ZN(n3478) );
  NAND2_X1 U3357 ( .A1(n1672), .A2(n1674), .ZN(n3479) );
  NAND2_X1 U3358 ( .A1(n1699), .A2(n1674), .ZN(n3480) );
  NAND3_X1 U3359 ( .A1(n3478), .A2(n3480), .A3(n3479), .ZN(n1669) );
  NOR2_X4 U3360 ( .A1(n3481), .A2(n3724), .ZN(n3751) );
  XNOR2_X1 U3361 ( .A(a[16]), .B(n345), .ZN(n3481) );
  NAND2_X4 U3362 ( .A1(n3690), .A2(n3691), .ZN(n3724) );
  NOR2_X1 U3363 ( .A1(n1842), .A2(n1861), .ZN(n864) );
  NAND2_X1 U3364 ( .A1(n3460), .A2(n851), .ZN(n842) );
  NAND2_X1 U3365 ( .A1(n1011), .A2(n815), .ZN(n565) );
  NAND2_X1 U3366 ( .A1(n1642), .A2(n1669), .ZN(n815) );
  INV_X1 U3367 ( .A(n1486), .ZN(n1487) );
  NOR2_X1 U3368 ( .A1(n2664), .A2(n3462), .ZN(n1486) );
  INV_X1 U3369 ( .A(n428), .ZN(n3482) );
  NAND2_X1 U3370 ( .A1(n998), .A2(n997), .ZN(n731) );
  OAI22_X1 U3371 ( .A1(n455), .A2(n2784), .B1(n2783), .B2(n3630), .ZN(n2214)
         );
  NOR2_X2 U3372 ( .A1(n1612), .A2(n1641), .ZN(n811) );
  OAI21_X1 U3373 ( .B1(n855), .B2(n849), .A(n850), .ZN(n848) );
  NAND2_X1 U3374 ( .A1(n851), .A2(n850), .ZN(n571) );
  INV_X1 U3375 ( .A(n850), .ZN(n852) );
  OAI22_X1 U3376 ( .A1(n455), .A2(n3730), .B1(n2799), .B2(n3630), .ZN(n2064)
         );
  XOR2_X1 U3377 ( .A(n2519), .B(n2487), .Z(n3483) );
  XOR2_X1 U3378 ( .A(n3483), .B(n2455), .Z(n1854) );
  NAND2_X1 U3379 ( .A1(n2455), .A2(n2519), .ZN(n3484) );
  NAND2_X1 U3380 ( .A1(n2455), .A2(n2487), .ZN(n3485) );
  NAND2_X1 U3381 ( .A1(n2519), .A2(n2487), .ZN(n3486) );
  NAND3_X1 U3382 ( .A1(n3484), .A2(n3486), .A3(n3485), .ZN(n1853) );
  OAI22_X1 U3383 ( .A1(n428), .A2(n3080), .B1(n3079), .B2(n3664), .ZN(n2519)
         );
  AOI21_X1 U3384 ( .B1(n786), .B2(n3618), .A(n787), .ZN(n3487) );
  XOR2_X1 U3385 ( .A(n1583), .B(n1555), .Z(n3488) );
  XOR2_X2 U3386 ( .A(n1553), .B(n3488), .Z(n1551) );
  NAND2_X1 U3387 ( .A1(n1553), .A2(n1583), .ZN(n3489) );
  NAND2_X1 U3388 ( .A1(n1553), .A2(n1555), .ZN(n3490) );
  NAND2_X1 U3389 ( .A1(n1583), .A2(n1555), .ZN(n3491) );
  NAND3_X1 U3390 ( .A1(n3489), .A2(n3491), .A3(n3490), .ZN(n1550) );
  AOI21_X1 U3391 ( .B1(n786), .B2(n799), .A(n787), .ZN(n785) );
  NAND2_X2 U3392 ( .A1(n1551), .A2(n1581), .ZN(n801) );
  INV_X1 U3393 ( .A(n840), .ZN(n838) );
  NAND2_X1 U3394 ( .A1(n3679), .A2(n840), .ZN(n569) );
  OAI22_X1 U3395 ( .A1(n3065), .A2(n428), .B1(n3064), .B2(n3664), .ZN(n2504)
         );
  BUF_X1 U3396 ( .A(n811), .Z(n3492) );
  NOR2_X1 U3397 ( .A1(n3445), .A2(n1641), .ZN(n3517) );
  BUF_X1 U3398 ( .A(n753), .Z(n3493) );
  NAND2_X1 U3399 ( .A1(n1351), .A2(n1376), .ZN(n760) );
  OAI22_X1 U3400 ( .A1(n419), .A2(n3165), .B1(n3164), .B2(n3511), .ZN(n2607)
         );
  INV_X2 U3401 ( .A(n3699), .ZN(n3700) );
  XNOR2_X1 U3402 ( .A(a[14]), .B(n342), .ZN(n3546) );
  XOR2_X1 U3403 ( .A(a[24]), .B(n357), .Z(n3231) );
  NAND2_X1 U3404 ( .A1(n757), .A2(n3446), .ZN(n555) );
  INV_X1 U3405 ( .A(n760), .ZN(n758) );
  NAND2_X1 U3406 ( .A1(n1010), .A2(n812), .ZN(n564) );
  XOR2_X1 U3407 ( .A(n1877), .B(n1879), .Z(n3494) );
  XOR2_X1 U3408 ( .A(n3494), .B(n1875), .Z(n1852) );
  XOR2_X1 U3409 ( .A(n1869), .B(n1867), .Z(n3495) );
  XOR2_X1 U3410 ( .A(n3495), .B(n1852), .Z(n1846) );
  NAND2_X1 U3411 ( .A1(n1877), .A2(n1879), .ZN(n3496) );
  NAND2_X1 U3412 ( .A1(n1877), .A2(n1875), .ZN(n3497) );
  NAND2_X1 U3413 ( .A1(n1879), .A2(n1875), .ZN(n3498) );
  NAND3_X1 U3414 ( .A1(n3496), .A2(n3497), .A3(n3498), .ZN(n1851) );
  NAND2_X1 U3415 ( .A1(n1869), .A2(n1867), .ZN(n3499) );
  NAND2_X1 U3416 ( .A1(n1869), .A2(n1852), .ZN(n3500) );
  NAND2_X1 U3417 ( .A1(n1867), .A2(n1852), .ZN(n3501) );
  NAND3_X1 U3418 ( .A1(n3499), .A2(n3500), .A3(n3501), .ZN(n1845) );
  OR2_X1 U3419 ( .A1(n3693), .A2(n3019), .ZN(n3502) );
  OR2_X1 U3420 ( .A1(n3018), .A2(n3566), .ZN(n3503) );
  NAND2_X1 U3421 ( .A1(n3502), .A2(n3503), .ZN(n2456) );
  INV_X2 U3422 ( .A(n3734), .ZN(n3693) );
  XNOR2_X1 U3423 ( .A(n489), .B(n336), .ZN(n3018) );
  XOR2_X1 U3424 ( .A(n1460), .B(n1435), .Z(n3504) );
  XOR2_X1 U3425 ( .A(n1433), .B(n3504), .Z(n1431) );
  NAND2_X1 U3426 ( .A1(n1433), .A2(n1460), .ZN(n3505) );
  NAND2_X1 U3427 ( .A1(n1433), .A2(n1435), .ZN(n3506) );
  NAND2_X1 U3428 ( .A1(n1460), .A2(n1435), .ZN(n3507) );
  NAND3_X1 U3429 ( .A1(n3505), .A2(n3507), .A3(n3506), .ZN(n1430) );
  INV_X1 U3430 ( .A(n3424), .ZN(n3508) );
  NAND2_X1 U3431 ( .A1(n1403), .A2(n1430), .ZN(n773) );
  NAND2_X1 U3432 ( .A1(n1003), .A2(n3473), .ZN(n557) );
  OAI22_X1 U3433 ( .A1(n455), .A2(n2776), .B1(n2775), .B2(n3630), .ZN(n2206)
         );
  NAND2_X2 U3434 ( .A1(n694), .A2(n994), .ZN(n692) );
  AOI21_X2 U3435 ( .B1(n694), .B2(n703), .A(n695), .ZN(n693) );
  AND2_X2 U3436 ( .A1(n1281), .A2(n1302), .ZN(n3509) );
  INV_X4 U3437 ( .A(n3509), .ZN(n739) );
  INV_X2 U3438 ( .A(n369), .ZN(n3510) );
  INV_X8 U3439 ( .A(n3510), .ZN(n3511) );
  NOR2_X2 U3440 ( .A1(n731), .A2(n747), .ZN(n729) );
  INV_X1 U3441 ( .A(n747), .ZN(n999) );
  NAND2_X1 U3442 ( .A1(n736), .A2(n997), .ZN(n551) );
  INV_X1 U3443 ( .A(n657), .ZN(n655) );
  OAI21_X1 U3444 ( .B1(n657), .B2(n637), .A(n638), .ZN(n636) );
  NOR2_X1 U3445 ( .A1(n1123), .A2(n1136), .ZN(n668) );
  NAND2_X2 U3446 ( .A1(n1123), .A2(n1136), .ZN(n669) );
  AOI21_X1 U3447 ( .B1(n876), .B2(n867), .A(n868), .ZN(n866) );
  NAND2_X2 U3448 ( .A1(n1303), .A2(n1326), .ZN(n748) );
  NOR2_X2 U3449 ( .A1(n1303), .A2(n1326), .ZN(n747) );
  NAND2_X1 U3450 ( .A1(n3613), .A2(n770), .ZN(n556) );
  OAI21_X1 U3451 ( .B1(n773), .B2(n3409), .A(n770), .ZN(n768) );
  NOR2_X1 U3452 ( .A1(n1431), .A2(n1458), .ZN(n3651) );
  OAI21_X2 U3453 ( .B1(n3651), .B2(n781), .A(n778), .ZN(n3628) );
  INV_X1 U3454 ( .A(n363), .ZN(n3278) );
  XOR2_X1 U3455 ( .A(n2482), .B(n2546), .Z(n3513) );
  XOR2_X1 U3456 ( .A(n2450), .B(n3513), .Z(n1740) );
  NAND2_X1 U3457 ( .A1(n2450), .A2(n2482), .ZN(n3514) );
  NAND2_X1 U3458 ( .A1(n2450), .A2(n2546), .ZN(n3515) );
  NAND2_X1 U3459 ( .A1(n2482), .A2(n2546), .ZN(n3516) );
  NAND3_X1 U3460 ( .A1(n3514), .A2(n3516), .A3(n3515), .ZN(n1739) );
  OR2_X1 U3461 ( .A1(n434), .A2(n3013), .ZN(n3518) );
  OR2_X1 U3462 ( .A1(n3012), .A2(n3567), .ZN(n3519) );
  NAND2_X1 U3463 ( .A1(n3518), .A2(n3519), .ZN(n2450) );
  OAI22_X1 U3464 ( .A1(n3602), .A2(n3044), .B1(n3043), .B2(n381), .ZN(n2482)
         );
  XNOR2_X1 U3465 ( .A(n499), .B(n336), .ZN(n3013) );
  XNOR2_X1 U3466 ( .A(n501), .B(n336), .ZN(n3012) );
  INV_X2 U3467 ( .A(n3564), .ZN(n3567) );
  OAI22_X1 U3468 ( .A1(n428), .A2(n3066), .B1(n3065), .B2(n3664), .ZN(n2505)
         );
  AOI21_X2 U3469 ( .B1(n3628), .B2(n767), .A(n768), .ZN(n766) );
  INV_X2 U3470 ( .A(n411), .ZN(n3520) );
  INV_X1 U3471 ( .A(n3520), .ZN(n3521) );
  INV_X2 U3472 ( .A(n3520), .ZN(n3523) );
  INV_X2 U3473 ( .A(n3520), .ZN(n3522) );
  INV_X1 U3474 ( .A(n690), .ZN(n688) );
  AOI21_X1 U3475 ( .B1(n3460), .B2(n852), .A(n845), .ZN(n3524) );
  INV_X1 U3476 ( .A(n419), .ZN(n3525) );
  INV_X2 U3477 ( .A(n3525), .ZN(n3526) );
  AOI21_X1 U3478 ( .B1(n3460), .B2(n852), .A(n845), .ZN(n843) );
  OAI22_X1 U3479 ( .A1(n419), .A2(n3164), .B1(n3163), .B2(n3511), .ZN(n2606)
         );
  NOR2_X1 U3480 ( .A1(n1219), .A2(n1238), .ZN(n715) );
  NAND2_X1 U3481 ( .A1(n1219), .A2(n1238), .ZN(n716) );
  NAND2_X2 U3482 ( .A1(n996), .A2(n995), .ZN(n711) );
  AND2_X1 U3483 ( .A1(n465), .A2(a[0]), .ZN(product[0]) );
  NAND2_X1 U3484 ( .A1(n1491), .A2(n1520), .ZN(n3527) );
  NAND2_X1 U3485 ( .A1(n1491), .A2(n1493), .ZN(n3528) );
  NAND2_X1 U3486 ( .A1(n1520), .A2(n1493), .ZN(n3529) );
  NAND3_X1 U3487 ( .A1(n3527), .A2(n3529), .A3(n3528), .ZN(n1488) );
  NAND2_X1 U3488 ( .A1(n998), .A2(n739), .ZN(n552) );
  BUF_X1 U3489 ( .A(n775), .Z(n3530) );
  INV_X1 U3490 ( .A(n3533), .ZN(n3531) );
  AND2_X1 U3491 ( .A1(n3677), .A2(n3678), .ZN(n3532) );
  AND2_X4 U3492 ( .A1(n3677), .A2(n3678), .ZN(n3533) );
  INV_X1 U3493 ( .A(n897), .ZN(n896) );
  NAND2_X1 U3494 ( .A1(n1964), .A2(n1977), .ZN(n908) );
  OAI21_X1 U3495 ( .B1(a[0]), .B2(n3589), .A(n321), .ZN(n2604) );
  NAND2_X1 U3496 ( .A1(n885), .A2(n888), .ZN(n577) );
  NAND2_X1 U3497 ( .A1(n885), .A2(n892), .ZN(n883) );
  AOI21_X2 U3498 ( .B1(n885), .B2(n893), .A(n886), .ZN(n884) );
  INV_X1 U3499 ( .A(n887), .ZN(n885) );
  INV_X1 U3500 ( .A(n738), .ZN(n998) );
  OAI22_X1 U3501 ( .A1(n3474), .A2(n2846), .B1(n2845), .B2(n3672), .ZN(n2278)
         );
  NOR2_X2 U3502 ( .A1(n800), .A2(n803), .ZN(n798) );
  OAI22_X1 U3503 ( .A1(n3601), .A2(n3048), .B1(n3047), .B2(n381), .ZN(n2486)
         );
  OAI22_X1 U3504 ( .A1(n3601), .A2(n3288), .B1(n3063), .B2(n381), .ZN(n2072)
         );
  OAI22_X1 U3505 ( .A1(n3601), .A2(n3059), .B1(n3058), .B2(n381), .ZN(n2497)
         );
  OAI22_X1 U3506 ( .A1(n3601), .A2(n3040), .B1(n3039), .B2(n381), .ZN(n2478)
         );
  OAI22_X1 U3507 ( .A1(n3601), .A2(n3045), .B1(n3044), .B2(n381), .ZN(n2483)
         );
  OAI22_X1 U3508 ( .A1(n3601), .A2(n3052), .B1(n3051), .B2(n381), .ZN(n2490)
         );
  OAI22_X1 U3509 ( .A1(n3601), .A2(n3049), .B1(n3048), .B2(n381), .ZN(n2487)
         );
  OAI22_X1 U3510 ( .A1(n3601), .A2(n3053), .B1(n3052), .B2(n381), .ZN(n2491)
         );
  OAI22_X1 U3511 ( .A1(n3601), .A2(n3035), .B1(n3034), .B2(n381), .ZN(n2473)
         );
  OAI22_X1 U3512 ( .A1(n3601), .A2(n3034), .B1(n3033), .B2(n381), .ZN(n2472)
         );
  NAND2_X4 U3513 ( .A1(n3688), .A2(n342), .ZN(n3691) );
  NOR2_X1 U3514 ( .A1(n2662), .A2(n3462), .ZN(n1428) );
  INV_X1 U3515 ( .A(n1428), .ZN(n1429) );
  XOR2_X1 U3516 ( .A(n2218), .B(n2410), .Z(n3534) );
  XOR2_X2 U3517 ( .A(n3534), .B(n2186), .Z(n1513) );
  XOR2_X1 U3518 ( .A(n1515), .B(n1511), .Z(n3535) );
  XOR2_X1 U3519 ( .A(n3535), .B(n1513), .Z(n1501) );
  NAND2_X1 U3520 ( .A1(n2218), .A2(n2410), .ZN(n3536) );
  NAND2_X1 U3521 ( .A1(n2218), .A2(n2186), .ZN(n3537) );
  NAND2_X1 U3522 ( .A1(n2410), .A2(n2186), .ZN(n3538) );
  NAND3_X1 U3523 ( .A1(n3536), .A2(n3537), .A3(n3538), .ZN(n1512) );
  NAND2_X1 U3524 ( .A1(n1515), .A2(n1511), .ZN(n3539) );
  NAND2_X1 U3525 ( .A1(n1515), .A2(n1513), .ZN(n3540) );
  NAND2_X1 U3526 ( .A1(n1511), .A2(n1513), .ZN(n3541) );
  NAND3_X1 U3527 ( .A1(n3539), .A2(n3540), .A3(n3541), .ZN(n1500) );
  OR2_X1 U3528 ( .A1(n455), .A2(n2788), .ZN(n3542) );
  OR2_X1 U3529 ( .A1(n2787), .A2(n3631), .ZN(n3543) );
  NAND2_X2 U3530 ( .A1(n3542), .A2(n3543), .ZN(n2218) );
  XNOR2_X1 U3531 ( .A(n489), .B(n357), .ZN(n2787) );
  INV_X4 U3532 ( .A(n3649), .ZN(n3631) );
  INV_X1 U3533 ( .A(n1003), .ZN(n3544) );
  INV_X1 U3534 ( .A(n3707), .ZN(n3545) );
  INV_X4 U3535 ( .A(n3734), .ZN(n3552) );
  NOR2_X2 U3536 ( .A1(n869), .A2(n874), .ZN(n867) );
  NOR2_X1 U3537 ( .A1(n1882), .A2(n1899), .ZN(n874) );
  INV_X1 U3538 ( .A(n3700), .ZN(n390) );
  OAI21_X1 U3539 ( .B1(n896), .B2(n883), .A(n884), .ZN(n882) );
  XNOR2_X2 U3540 ( .A(n3512), .B(n3745), .ZN(n3547) );
  INV_X4 U3541 ( .A(n3547), .ZN(n3744) );
  AOI21_X1 U3542 ( .B1(n603), .B2(n980), .A(n600), .ZN(n598) );
  OAI22_X1 U3543 ( .A1(n3720), .A2(n2726), .B1(n2725), .B2(n3522), .ZN(n2154)
         );
  OAI22_X1 U3544 ( .A1(n3720), .A2(n2732), .B1(n2731), .B2(n3523), .ZN(n2160)
         );
  OAI22_X1 U3545 ( .A1(n3720), .A2(n3278), .B1(n2733), .B2(n3523), .ZN(n2062)
         );
  OAI22_X1 U3546 ( .A1(n3720), .A2(n2716), .B1(n2715), .B2(n3522), .ZN(n2144)
         );
  OAI22_X1 U3547 ( .A1(n3720), .A2(n2727), .B1(n2726), .B2(n3522), .ZN(n2155)
         );
  INV_X4 U3548 ( .A(n3706), .ZN(n411) );
  INV_X1 U3549 ( .A(n819), .ZN(n1012) );
  AOI21_X1 U3550 ( .B1(n826), .B2(n817), .A(n818), .ZN(n816) );
  AOI21_X1 U3551 ( .B1(n809), .B2(n818), .A(n810), .ZN(n808) );
  XNOR2_X1 U3552 ( .A(n3732), .B(n3548), .ZN(product[62]) );
  AND2_X1 U3553 ( .A1(n979), .A2(n597), .ZN(n3548) );
  AND2_X2 U3554 ( .A1(n3243), .A2(n3511), .ZN(n3589) );
  XOR2_X1 U3555 ( .A(a[0]), .B(n321), .Z(n3243) );
  OAI21_X1 U3556 ( .B1(n604), .B2(n531), .A(n605), .ZN(n3704) );
  INV_X2 U3557 ( .A(n3652), .ZN(n3655) );
  BUF_X1 U3558 ( .A(n801), .Z(n3549) );
  INV_X4 U3559 ( .A(n3734), .ZN(n3551) );
  AND2_X4 U3560 ( .A1(n3238), .A2(n3565), .ZN(n3734) );
  OAI21_X1 U3561 ( .B1(n3608), .B2(n750), .A(n751), .ZN(n3555) );
  NOR2_X2 U3562 ( .A1(n1551), .A2(n1581), .ZN(n3556) );
  OAI21_X1 U3563 ( .B1(n3608), .B2(n750), .A(n751), .ZN(n749) );
  NOR2_X1 U3564 ( .A1(n1551), .A2(n1581), .ZN(n800) );
  INV_X1 U3565 ( .A(n3608), .ZN(n3557) );
  INV_X2 U3566 ( .A(n3558), .ZN(n3559) );
  AOI21_X2 U3567 ( .B1(n859), .B2(n868), .A(n860), .ZN(n858) );
  OAI22_X1 U3568 ( .A1(n3471), .A2(n2797), .B1(n2796), .B2(n3630), .ZN(n2227)
         );
  NOR2_X2 U3569 ( .A1(n1670), .A2(n1697), .ZN(n819) );
  NOR2_X2 U3570 ( .A1(n814), .A2(n3517), .ZN(n809) );
  AOI21_X1 U3571 ( .B1(n3555), .B2(n999), .A(n746), .ZN(n3560) );
  BUF_X1 U3572 ( .A(n829), .Z(n3561) );
  AOI21_X1 U3573 ( .B1(n749), .B2(n999), .A(n746), .ZN(n744) );
  BUF_X1 U3574 ( .A(n780), .Z(n3562) );
  NOR2_X1 U3575 ( .A1(n1488), .A2(n1459), .ZN(n780) );
  XNOR2_X1 U3576 ( .A(n1554), .B(n3563), .ZN(n1521) );
  XNOR2_X1 U3577 ( .A(n1525), .B(n1556), .ZN(n3563) );
  OAI22_X1 U3578 ( .A1(n446), .A2(n2888), .B1(n2887), .B2(n396), .ZN(n2321) );
  NOR2_X2 U3579 ( .A1(n1820), .A2(n1841), .ZN(n861) );
  OAI22_X1 U3580 ( .A1(n443), .A2(n2907), .B1(n2906), .B2(n393), .ZN(n2341) );
  OAI22_X1 U3581 ( .A1(n443), .A2(n2904), .B1(n2903), .B2(n393), .ZN(n2338) );
  OAI22_X1 U3582 ( .A1(n443), .A2(n2925), .B1(n2924), .B2(n393), .ZN(n2359) );
  OAI22_X1 U3583 ( .A1(n443), .A2(n2905), .B1(n2904), .B2(n393), .ZN(n2339) );
  OAI22_X1 U3584 ( .A1(n443), .A2(n2906), .B1(n2905), .B2(n393), .ZN(n2340) );
  OAI22_X1 U3585 ( .A1(n443), .A2(n2917), .B1(n2916), .B2(n393), .ZN(n2351) );
  OAI22_X1 U3586 ( .A1(n3623), .A2(n2927), .B1(n2926), .B2(n393), .ZN(n2361)
         );
  OAI22_X1 U3587 ( .A1(n3623), .A2(n2916), .B1(n2915), .B2(n393), .ZN(n2350)
         );
  OAI22_X1 U3588 ( .A1(n443), .A2(n2912), .B1(n2911), .B2(n393), .ZN(n2346) );
  OAI22_X1 U3589 ( .A1(n443), .A2(n2915), .B1(n2914), .B2(n393), .ZN(n2349) );
  OAI22_X1 U3590 ( .A1(n3623), .A2(n2910), .B1(n2909), .B2(n393), .ZN(n2344)
         );
  OAI22_X1 U3591 ( .A1(n3623), .A2(n2922), .B1(n2921), .B2(n393), .ZN(n2356)
         );
  OAI22_X1 U3592 ( .A1(n443), .A2(n2921), .B1(n2920), .B2(n393), .ZN(n2355) );
  OAI22_X1 U3593 ( .A1(n3623), .A2(n2911), .B1(n2910), .B2(n393), .ZN(n2345)
         );
  OAI22_X1 U3594 ( .A1(n3623), .A2(n2899), .B1(n393), .B2(n3416), .ZN(n2333)
         );
  OAI22_X1 U3595 ( .A1(n3623), .A2(n2908), .B1(n2907), .B2(n393), .ZN(n2342)
         );
  AOI21_X2 U3596 ( .B1(n3710), .B2(n654), .A(n655), .ZN(n3726) );
  NOR2_X2 U3597 ( .A1(n1519), .A2(n1550), .ZN(n793) );
  INV_X2 U3598 ( .A(n384), .ZN(n3564) );
  INV_X1 U3599 ( .A(n3564), .ZN(n3565) );
  INV_X2 U3600 ( .A(n3564), .ZN(n3566) );
  NAND2_X1 U3601 ( .A1(n1554), .A2(n1525), .ZN(n3568) );
  NAND2_X1 U3602 ( .A1(n1554), .A2(n1556), .ZN(n3569) );
  NAND2_X1 U3603 ( .A1(n1525), .A2(n1556), .ZN(n3570) );
  NAND3_X1 U3604 ( .A1(n3568), .A2(n3570), .A3(n3569), .ZN(n1520) );
  INV_X8 U3605 ( .A(n3738), .ZN(n3571) );
  INV_X1 U3606 ( .A(n3738), .ZN(n387) );
  INV_X8 U3607 ( .A(n3680), .ZN(n3667) );
  XOR2_X1 U3608 ( .A(a[12]), .B(n339), .Z(n3237) );
  INV_X1 U3609 ( .A(n3574), .ZN(n3572) );
  INV_X2 U3610 ( .A(n360), .ZN(n3279) );
  INV_X2 U3611 ( .A(n342), .ZN(n3689) );
  INV_X1 U3612 ( .A(n1009), .ZN(n3575) );
  INV_X1 U3613 ( .A(n3562), .ZN(n1005) );
  OAI22_X1 U3614 ( .A1(n3596), .A2(n3121), .B1(n3120), .B2(n3533), .ZN(n2561)
         );
  OAI22_X1 U3615 ( .A1(n3596), .A2(n3116), .B1(n3115), .B2(n3533), .ZN(n2556)
         );
  OAI22_X1 U3616 ( .A1(n3596), .A2(n3128), .B1(n3127), .B2(n3533), .ZN(n2568)
         );
  OAI22_X1 U3617 ( .A1(n3596), .A2(n3290), .B1(n3129), .B2(n3533), .ZN(n2074)
         );
  OAI22_X1 U3618 ( .A1(n3596), .A2(n3127), .B1(n3126), .B2(n3533), .ZN(n2567)
         );
  OAI22_X1 U3619 ( .A1(n3596), .A2(n3125), .B1(n3124), .B2(n3533), .ZN(n2565)
         );
  OAI22_X1 U3620 ( .A1(n3596), .A2(n3126), .B1(n3125), .B2(n3533), .ZN(n2566)
         );
  OAI22_X1 U3621 ( .A1(n3596), .A2(n3123), .B1(n3122), .B2(n3533), .ZN(n2563)
         );
  OAI22_X1 U3622 ( .A1(n3596), .A2(n3119), .B1(n3118), .B2(n3533), .ZN(n2559)
         );
  OAI22_X1 U3623 ( .A1(n3596), .A2(n3124), .B1(n3123), .B2(n3533), .ZN(n2564)
         );
  OAI22_X1 U3624 ( .A1(n3596), .A2(n3108), .B1(n3107), .B2(n3533), .ZN(n2548)
         );
  OAI22_X1 U3625 ( .A1(n3596), .A2(n3122), .B1(n3121), .B2(n3533), .ZN(n2562)
         );
  OAI22_X1 U3626 ( .A1(n3596), .A2(n3117), .B1(n3116), .B2(n3533), .ZN(n2557)
         );
  OAI22_X1 U3627 ( .A1(n3596), .A2(n3114), .B1(n3113), .B2(n3533), .ZN(n2554)
         );
  OAI22_X1 U3628 ( .A1(n3596), .A2(n3120), .B1(n3119), .B2(n3533), .ZN(n2560)
         );
  OAI22_X1 U3629 ( .A1(n3596), .A2(n3105), .B1(n3104), .B2(n3533), .ZN(n2545)
         );
  OAI22_X1 U3630 ( .A1(n3596), .A2(n3109), .B1(n3108), .B2(n3533), .ZN(n2549)
         );
  OAI22_X1 U3631 ( .A1(n3596), .A2(n3112), .B1(n3111), .B2(n3533), .ZN(n2552)
         );
  OAI22_X1 U3632 ( .A1(n3596), .A2(n3113), .B1(n3112), .B2(n3533), .ZN(n2553)
         );
  OAI22_X1 U3633 ( .A1(n3596), .A2(n3103), .B1(n3102), .B2(n3533), .ZN(n2543)
         );
  OAI22_X1 U3634 ( .A1(n3596), .A2(n3110), .B1(n3109), .B2(n3533), .ZN(n2550)
         );
  OAI22_X1 U3635 ( .A1(n3596), .A2(n3111), .B1(n3110), .B2(n3533), .ZN(n2551)
         );
  OAI22_X1 U3636 ( .A1(n3596), .A2(n3104), .B1(n3103), .B2(n3533), .ZN(n2544)
         );
  OAI22_X1 U3637 ( .A1(n3596), .A2(n3102), .B1(n3101), .B2(n3533), .ZN(n2542)
         );
  OAI22_X1 U3638 ( .A1(n3596), .A2(n3101), .B1(n3100), .B2(n3533), .ZN(n2541)
         );
  OAI22_X1 U3639 ( .A1(n3596), .A2(n3106), .B1(n3105), .B2(n3533), .ZN(n2546)
         );
  OAI22_X1 U3640 ( .A1(n3596), .A2(n3118), .B1(n3117), .B2(n3533), .ZN(n2558)
         );
  OAI22_X1 U3641 ( .A1(n3596), .A2(n3107), .B1(n3106), .B2(n3533), .ZN(n2547)
         );
  OAI22_X1 U3642 ( .A1(n3596), .A2(n3115), .B1(n3114), .B2(n3533), .ZN(n2555)
         );
  OAI22_X1 U3643 ( .A1(n3596), .A2(n3099), .B1(n3098), .B2(n3533), .ZN(n2539)
         );
  AND2_X2 U3644 ( .A1(n3424), .A2(n3577), .ZN(n3576) );
  INV_X8 U3645 ( .A(n3576), .ZN(n428) );
  XOR2_X1 U3646 ( .A(n2348), .B(n2124), .Z(n3578) );
  XOR2_X2 U3647 ( .A(n3578), .B(n2188), .Z(n1577) );
  XOR2_X1 U3648 ( .A(n1571), .B(n1573), .Z(n3579) );
  XOR2_X1 U3649 ( .A(n3579), .B(n1577), .Z(n1563) );
  NAND2_X1 U3650 ( .A1(n2348), .A2(n2124), .ZN(n3580) );
  NAND2_X1 U3651 ( .A1(n2348), .A2(n2188), .ZN(n3581) );
  NAND2_X1 U3652 ( .A1(n3586), .A2(n2188), .ZN(n3582) );
  NAND3_X1 U3653 ( .A1(n3580), .A2(n3581), .A3(n3582), .ZN(n1576) );
  NAND2_X1 U3654 ( .A1(n1571), .A2(n1573), .ZN(n3583) );
  NAND2_X1 U3655 ( .A1(n1571), .A2(n1577), .ZN(n3584) );
  NAND2_X1 U3656 ( .A1(n1573), .A2(n1577), .ZN(n3585) );
  NAND3_X1 U3657 ( .A1(n3583), .A2(n3584), .A3(n3585), .ZN(n1562) );
  BUF_X1 U3658 ( .A(n2124), .Z(n3586) );
  INV_X1 U3659 ( .A(n803), .ZN(n1009) );
  AND2_X2 U3660 ( .A1(n3588), .A2(n399), .ZN(n3587) );
  INV_X2 U3661 ( .A(n399), .ZN(n3671) );
  INV_X8 U3662 ( .A(n3589), .ZN(n419) );
  OAI22_X1 U3663 ( .A1(n419), .A2(n3166), .B1(n3165), .B2(n3511), .ZN(n2608)
         );
  OAI22_X1 U3664 ( .A1(n464), .A2(n2673), .B1(n2672), .B2(n3654), .ZN(n2100)
         );
  OAI22_X1 U3665 ( .A1(n464), .A2(n2675), .B1(n2674), .B2(n3655), .ZN(n2102)
         );
  OAI22_X1 U3666 ( .A1(n464), .A2(n2681), .B1(n2680), .B2(n3654), .ZN(n2108)
         );
  OAI22_X1 U3667 ( .A1(n464), .A2(n2676), .B1(n2675), .B2(n3655), .ZN(n2103)
         );
  OAI22_X1 U3668 ( .A1(n464), .A2(n2690), .B1(n2689), .B2(n3654), .ZN(n2117)
         );
  OAI22_X1 U3669 ( .A1(n464), .A2(n2680), .B1(n2679), .B2(n3654), .ZN(n2107)
         );
  OAI22_X1 U3670 ( .A1(n464), .A2(n2679), .B1(n2678), .B2(n3655), .ZN(n2106)
         );
  OAI22_X1 U3671 ( .A1(n464), .A2(n2689), .B1(n2688), .B2(n3654), .ZN(n2116)
         );
  OAI22_X1 U3672 ( .A1(n464), .A2(n2688), .B1(n2687), .B2(n3654), .ZN(n2115)
         );
  OAI22_X1 U3673 ( .A1(n464), .A2(n2686), .B1(n2685), .B2(n3655), .ZN(n2113)
         );
  OAI22_X1 U3674 ( .A1(n464), .A2(n2678), .B1(n2677), .B2(n3655), .ZN(n2105)
         );
  OAI22_X1 U3675 ( .A1(n464), .A2(n2684), .B1(n2683), .B2(n3654), .ZN(n2111)
         );
  OAI22_X1 U3676 ( .A1(n464), .A2(n2683), .B1(n2682), .B2(n3655), .ZN(n2110)
         );
  OAI22_X1 U3677 ( .A1(n464), .A2(n2695), .B1(n2694), .B2(n3655), .ZN(n2122)
         );
  OAI22_X1 U3678 ( .A1(n464), .A2(n2692), .B1(n2691), .B2(n3654), .ZN(n2119)
         );
  OAI22_X1 U3679 ( .A1(n464), .A2(n2677), .B1(n2676), .B2(n3654), .ZN(n2104)
         );
  OAI22_X1 U3680 ( .A1(n464), .A2(n2687), .B1(n2686), .B2(n3655), .ZN(n2114)
         );
  OAI22_X1 U3681 ( .A1(n464), .A2(n2694), .B1(n2693), .B2(n3655), .ZN(n2121)
         );
  OAI22_X1 U3682 ( .A1(n464), .A2(n2685), .B1(n2684), .B2(n3655), .ZN(n2112)
         );
  OAI22_X1 U3683 ( .A1(n464), .A2(n2682), .B1(n2681), .B2(n3654), .ZN(n2109)
         );
  OAI22_X1 U3684 ( .A1(n464), .A2(n2693), .B1(n2692), .B2(n3654), .ZN(n2120)
         );
  OAI22_X1 U3685 ( .A1(n464), .A2(n2691), .B1(n2690), .B2(n3655), .ZN(n2118)
         );
  OAI22_X1 U3686 ( .A1(n464), .A2(n2698), .B1(n2697), .B2(n3654), .ZN(n2125)
         );
  OAI22_X1 U3687 ( .A1(n464), .A2(n2696), .B1(n2695), .B2(n3654), .ZN(n2123)
         );
  OAI22_X1 U3688 ( .A1(n464), .A2(n2697), .B1(n2696), .B2(n3655), .ZN(n2124)
         );
  OAI22_X1 U3689 ( .A1(n464), .A2(n3462), .B1(n2700), .B2(n3654), .ZN(n2061)
         );
  OAI22_X1 U3690 ( .A1(n3667), .A2(n2976), .B1(n2975), .B2(n3571), .ZN(n2412)
         );
  INV_X1 U3691 ( .A(n3493), .ZN(n751) );
  NOR2_X2 U3692 ( .A1(n754), .A2(n759), .ZN(n752) );
  OAI22_X1 U3693 ( .A1(n461), .A2(n2701), .B1(n3523), .B2(n3278), .ZN(n2129)
         );
  OAI22_X1 U3694 ( .A1(n461), .A2(n2703), .B1(n2702), .B2(n3522), .ZN(n2131)
         );
  OAI22_X1 U3695 ( .A1(n461), .A2(n2704), .B1(n2703), .B2(n3522), .ZN(n2132)
         );
  OAI22_X1 U3696 ( .A1(n461), .A2(n2706), .B1(n2705), .B2(n3522), .ZN(n2134)
         );
  OAI22_X1 U3697 ( .A1(n461), .A2(n2712), .B1(n2711), .B2(n3522), .ZN(n2140)
         );
  OAI22_X1 U3698 ( .A1(n461), .A2(n2707), .B1(n2706), .B2(n3522), .ZN(n2135)
         );
  OAI22_X1 U3699 ( .A1(n461), .A2(n2711), .B1(n2710), .B2(n3523), .ZN(n2139)
         );
  OAI22_X1 U3700 ( .A1(n461), .A2(n2718), .B1(n2717), .B2(n3522), .ZN(n2146)
         );
  OAI22_X1 U3701 ( .A1(n461), .A2(n2715), .B1(n2714), .B2(n3523), .ZN(n2143)
         );
  OAI22_X1 U3702 ( .A1(n461), .A2(n2714), .B1(n2713), .B2(n3522), .ZN(n2142)
         );
  OAI22_X1 U3703 ( .A1(n461), .A2(n2723), .B1(n2722), .B2(n3523), .ZN(n2151)
         );
  XOR2_X1 U3704 ( .A(n1775), .B(n1754), .Z(n3590) );
  XOR2_X1 U3705 ( .A(n1752), .B(n3590), .Z(n1750) );
  NAND2_X1 U3706 ( .A1(n1752), .A2(n1775), .ZN(n3591) );
  NAND2_X1 U3707 ( .A1(n1752), .A2(n1754), .ZN(n3592) );
  NAND2_X1 U3708 ( .A1(n1775), .A2(n1754), .ZN(n3593) );
  NAND3_X1 U3709 ( .A1(n3591), .A2(n3593), .A3(n3592), .ZN(n1749) );
  OR2_X2 U3710 ( .A1(n1750), .A2(n1773), .ZN(n3679) );
  NAND2_X1 U3711 ( .A1(n1750), .A2(n1773), .ZN(n840) );
  INV_X1 U3712 ( .A(n3705), .ZN(n3594) );
  INV_X4 U3713 ( .A(n3748), .ZN(n3595) );
  AND2_X4 U3714 ( .A1(n3230), .A2(n3594), .ZN(n3748) );
  INV_X4 U3715 ( .A(n3695), .ZN(n384) );
  OAI21_X2 U3716 ( .B1(n754), .B2(n760), .A(n755), .ZN(n753) );
  NOR2_X2 U3717 ( .A1(n1327), .A2(n1350), .ZN(n754) );
  OAI22_X1 U3718 ( .A1(n428), .A2(n3064), .B1(n3664), .B2(n3289), .ZN(n2503)
         );
  INV_X8 U3719 ( .A(n3724), .ZN(n393) );
  INV_X8 U3720 ( .A(n3684), .ZN(n3596) );
  INV_X1 U3721 ( .A(n3684), .ZN(n425) );
  INV_X1 U3722 ( .A(n735), .ZN(n997) );
  OAI22_X1 U3723 ( .A1(n434), .A2(n3016), .B1(n3015), .B2(n3567), .ZN(n2453)
         );
  OAI22_X1 U3724 ( .A1(n3552), .A2(n2999), .B1(n2998), .B2(n3567), .ZN(n2436)
         );
  OAI22_X1 U3725 ( .A1(n3552), .A2(n3011), .B1(n3010), .B2(n3567), .ZN(n2448)
         );
  OAI22_X1 U3726 ( .A1(n434), .A2(n3000), .B1(n2999), .B2(n3566), .ZN(n2437)
         );
  OAI22_X1 U3727 ( .A1(n3552), .A2(n3028), .B1(n3027), .B2(n3566), .ZN(n2465)
         );
  OAI22_X1 U3728 ( .A1(n3551), .A2(n3020), .B1(n3019), .B2(n3567), .ZN(n2457)
         );
  OAI22_X1 U3729 ( .A1(n434), .A2(n3014), .B1(n3013), .B2(n3567), .ZN(n2451)
         );
  OAI22_X1 U3730 ( .A1(n434), .A2(n3027), .B1(n3026), .B2(n3566), .ZN(n2464)
         );
  OAI22_X1 U3731 ( .A1(n3552), .A2(n3004), .B1(n3003), .B2(n3566), .ZN(n2441)
         );
  OAI22_X1 U3732 ( .A1(n3551), .A2(n3015), .B1(n3014), .B2(n3567), .ZN(n2452)
         );
  OAI22_X1 U3733 ( .A1(n3552), .A2(n3007), .B1(n3006), .B2(n3566), .ZN(n2444)
         );
  OAI22_X1 U3734 ( .A1(n434), .A2(n3001), .B1(n3000), .B2(n3566), .ZN(n2438)
         );
  INV_X2 U3735 ( .A(n390), .ZN(n3697) );
  NAND2_X1 U3736 ( .A1(n3420), .A2(n3597), .ZN(n3599) );
  NAND2_X1 U3737 ( .A1(n3598), .A2(n3599), .ZN(n3648) );
  INV_X1 U3738 ( .A(n3648), .ZN(n3681) );
  BUF_X1 U3739 ( .A(n3557), .Z(n3600) );
  NAND2_X2 U3740 ( .A1(n3239), .A2(n381), .ZN(n3602) );
  NAND2_X2 U3741 ( .A1(n3239), .A2(n381), .ZN(n3601) );
  INV_X1 U3742 ( .A(n3459), .ZN(n3743) );
  OAI22_X1 U3743 ( .A1(n3729), .A2(n2734), .B1(n408), .B2(n3572), .ZN(n2163)
         );
  OAI22_X1 U3744 ( .A1(n3693), .A2(n3005), .B1(n3004), .B2(n3567), .ZN(n2442)
         );
  BUF_X1 U3745 ( .A(n3555), .Z(n3603) );
  NAND2_X1 U3746 ( .A1(a[28]), .A2(n3279), .ZN(n3605) );
  NAND2_X2 U3747 ( .A1(n1934), .A2(n1949), .ZN(n891) );
  NOR2_X2 U3748 ( .A1(n1934), .A2(n1949), .ZN(n890) );
  INV_X1 U3749 ( .A(n339), .ZN(n3646) );
  NOR2_X2 U3750 ( .A1(n1642), .A2(n1669), .ZN(n814) );
  OAI22_X1 U3751 ( .A1(n3720), .A2(n2731), .B1(n2730), .B2(n3523), .ZN(n2159)
         );
  INV_X16 U3752 ( .A(n465), .ZN(n3752) );
  OAI21_X1 U3753 ( .B1(n866), .B2(n864), .A(n865), .ZN(n863) );
  INV_X1 U3754 ( .A(n864), .ZN(n1019) );
  NAND2_X2 U3755 ( .A1(n1842), .A2(n1861), .ZN(n865) );
  NAND2_X1 U3756 ( .A1(n1774), .A2(n1797), .ZN(n847) );
  OAI22_X1 U3757 ( .A1(n443), .A2(n2900), .B1(n2899), .B2(n393), .ZN(n2334) );
  OAI22_X1 U3758 ( .A1(n443), .A2(n2930), .B1(n2929), .B2(n393), .ZN(n2364) );
  OAI22_X1 U3759 ( .A1(n443), .A2(n3416), .B1(n2931), .B2(n393), .ZN(n2068) );
  OAI22_X1 U3760 ( .A1(n443), .A2(n2902), .B1(n2901), .B2(n393), .ZN(n2336) );
  OAI22_X1 U3761 ( .A1(n443), .A2(n2901), .B1(n2900), .B2(n393), .ZN(n2335) );
  OAI22_X1 U3762 ( .A1(n443), .A2(n2903), .B1(n2902), .B2(n393), .ZN(n2337) );
  OAI22_X1 U3763 ( .A1(n443), .A2(n2913), .B1(n2912), .B2(n393), .ZN(n2347) );
  OAI22_X1 U3764 ( .A1(n443), .A2(n2928), .B1(n2927), .B2(n393), .ZN(n2362) );
  OAI22_X1 U3765 ( .A1(n3623), .A2(n2918), .B1(n2917), .B2(n393), .ZN(n2352)
         );
  OAI22_X1 U3766 ( .A1(n3623), .A2(n2919), .B1(n2918), .B2(n393), .ZN(n2353)
         );
  OAI22_X1 U3767 ( .A1(n443), .A2(n2923), .B1(n2922), .B2(n393), .ZN(n2357) );
  OAI22_X1 U3768 ( .A1(n443), .A2(n2920), .B1(n2919), .B2(n393), .ZN(n2354) );
  OAI22_X1 U3769 ( .A1(n443), .A2(n2924), .B1(n2923), .B2(n393), .ZN(n2358) );
  OAI22_X1 U3770 ( .A1(n443), .A2(n2926), .B1(n2925), .B2(n393), .ZN(n2360) );
  OAI22_X1 U3771 ( .A1(n3623), .A2(n2909), .B1(n2908), .B2(n393), .ZN(n2343)
         );
  OAI22_X1 U3772 ( .A1(n3623), .A2(n2929), .B1(n2928), .B2(n393), .ZN(n2363)
         );
  AND2_X2 U3773 ( .A1(n3727), .A2(n3728), .ZN(n3608) );
  AND2_X2 U3774 ( .A1(n3727), .A2(n3728), .ZN(n531) );
  NAND2_X1 U3775 ( .A1(n1726), .A2(n1751), .ZN(n3609) );
  NAND2_X1 U3776 ( .A1(n1726), .A2(n1728), .ZN(n3610) );
  NAND2_X1 U3777 ( .A1(n1751), .A2(n1728), .ZN(n3611) );
  NAND3_X1 U3778 ( .A1(n3609), .A2(n3611), .A3(n3610), .ZN(n1723) );
  AOI21_X1 U3779 ( .B1(n828), .B2(n3442), .A(n3561), .ZN(n3612) );
  NAND2_X2 U3780 ( .A1(n1698), .A2(n1723), .ZN(n825) );
  NOR2_X1 U3781 ( .A1(n1698), .A2(n1723), .ZN(n824) );
  OR2_X2 U3782 ( .A1(n1724), .A2(n1749), .ZN(n3665) );
  AOI21_X1 U3783 ( .B1(n856), .B2(n828), .A(n829), .ZN(n827) );
  INV_X1 U3784 ( .A(n3410), .ZN(n1011) );
  OAI21_X1 U3785 ( .B1(n816), .B2(n3410), .A(n815), .ZN(n813) );
  OR2_X1 U3786 ( .A1(n1377), .A2(n1402), .ZN(n3613) );
  NAND2_X2 U3787 ( .A1(n3614), .A2(n351), .ZN(n3617) );
  NAND2_X2 U3788 ( .A1(n3616), .A2(n3617), .ZN(n3707) );
  OAI21_X1 U3789 ( .B1(n855), .B2(n842), .A(n3524), .ZN(n841) );
  OAI22_X1 U3790 ( .A1(n3458), .A2(n2954), .B1(n2953), .B2(n3698), .ZN(n2389)
         );
  OAI22_X1 U3791 ( .A1(n464), .A2(n2699), .B1(n2698), .B2(n3655), .ZN(n2126)
         );
  INV_X8 U3792 ( .A(n3685), .ZN(n464) );
  OAI21_X1 U3793 ( .B1(n3556), .B2(n804), .A(n801), .ZN(n3618) );
  NAND2_X2 U3794 ( .A1(n1582), .A2(n1611), .ZN(n804) );
  OAI22_X1 U3795 ( .A1(n3474), .A2(n2852), .B1(n2851), .B2(n3673), .ZN(n2284)
         );
  NOR2_X1 U3796 ( .A1(n1582), .A2(n1611), .ZN(n803) );
  NOR2_X2 U3797 ( .A1(n1281), .A2(n1302), .ZN(n738) );
  NAND2_X1 U3798 ( .A1(n3619), .A2(n3620), .ZN(n3622) );
  NAND2_X2 U3799 ( .A1(n3621), .A2(n3622), .ZN(n3738) );
  INV_X1 U3800 ( .A(n3739), .ZN(n3619) );
  INV_X1 U3801 ( .A(n336), .ZN(n3620) );
  INV_X4 U3802 ( .A(n3751), .ZN(n3623) );
  NAND2_X1 U3803 ( .A1(a[16]), .A2(n3689), .ZN(n3690) );
  NOR2_X1 U3804 ( .A1(n1351), .A2(n1376), .ZN(n759) );
  OAI21_X1 U3805 ( .B1(n728), .B2(n688), .A(n689), .ZN(n687) );
  NAND2_X1 U3806 ( .A1(n1327), .A2(n1350), .ZN(n755) );
  NAND2_X1 U3807 ( .A1(n3625), .A2(a[10]), .ZN(n3626) );
  NAND2_X1 U3808 ( .A1(n3624), .A2(n333), .ZN(n3627) );
  NAND2_X1 U3809 ( .A1(n3626), .A2(n3627), .ZN(n3719) );
  INV_X2 U3810 ( .A(n333), .ZN(n3625) );
  NAND2_X1 U3811 ( .A1(n859), .A2(n867), .ZN(n857) );
  NAND2_X1 U3812 ( .A1(n3665), .A2(n3679), .ZN(n830) );
  AOI21_X2 U3813 ( .B1(n3665), .B2(n838), .A(n833), .ZN(n831) );
  BUF_X1 U3814 ( .A(n781), .Z(n3629) );
  INV_X4 U3815 ( .A(n3649), .ZN(n3630) );
  NAND2_X1 U3816 ( .A1(n3472), .A2(n354), .ZN(n3634) );
  NAND2_X1 U3817 ( .A1(n3632), .A2(n3633), .ZN(n3635) );
  NAND2_X1 U3818 ( .A1(n3634), .A2(n3635), .ZN(n3735) );
  INV_X1 U3819 ( .A(n3472), .ZN(n3632) );
  INV_X1 U3820 ( .A(n3649), .ZN(n3650) );
  INV_X1 U3821 ( .A(n3735), .ZN(n405) );
  NAND2_X1 U3822 ( .A1(n3657), .A2(n357), .ZN(n3638) );
  NAND2_X1 U3823 ( .A1(n3636), .A2(n3637), .ZN(n3639) );
  NAND2_X2 U3824 ( .A1(n3638), .A2(n3639), .ZN(n3705) );
  INV_X1 U3825 ( .A(n3657), .ZN(n3636) );
  INV_X1 U3826 ( .A(n357), .ZN(n3637) );
  INV_X1 U3827 ( .A(n3522), .ZN(n3640) );
  OAI21_X1 U3828 ( .B1(n3608), .B2(n671), .A(n672), .ZN(n3641) );
  NAND2_X1 U3829 ( .A1(a[14]), .A2(n3643), .ZN(n3644) );
  NAND2_X1 U3830 ( .A1(n3642), .A2(n339), .ZN(n3645) );
  NAND2_X1 U3831 ( .A1(n3644), .A2(n3645), .ZN(n3725) );
  INV_X1 U3832 ( .A(a[14]), .ZN(n3642) );
  INV_X2 U3833 ( .A(n339), .ZN(n3643) );
  INV_X2 U3834 ( .A(n3646), .ZN(n3647) );
  INV_X2 U3835 ( .A(n3750), .ZN(n3670) );
  INV_X2 U3836 ( .A(n405), .ZN(n3649) );
  NOR2_X1 U3837 ( .A1(n1431), .A2(n1458), .ZN(n777) );
  NAND2_X1 U3838 ( .A1(n905), .A2(n900), .ZN(n898) );
  AOI21_X2 U3839 ( .B1(n906), .B2(n900), .A(n901), .ZN(n899) );
  OAI22_X1 U3840 ( .A1(n455), .A2(n2796), .B1(n2795), .B2(n3631), .ZN(n2226)
         );
  OAI21_X1 U3841 ( .B1(n843), .B2(n830), .A(n831), .ZN(n829) );
  NAND2_X1 U3842 ( .A1(n3708), .A2(n3549), .ZN(n562) );
  INV_X2 U3843 ( .A(n3547), .ZN(n3652) );
  INV_X1 U3844 ( .A(n3652), .ZN(n3653) );
  INV_X4 U3845 ( .A(n3652), .ZN(n3654) );
  NAND2_X1 U3846 ( .A1(n1519), .A2(n1550), .ZN(n794) );
  OAI22_X1 U3847 ( .A1(n3713), .A2(n2816), .B1(n2815), .B2(n402), .ZN(n2247)
         );
  OAI22_X1 U3848 ( .A1(n3713), .A2(n2804), .B1(n2803), .B2(n402), .ZN(n2235)
         );
  OAI22_X1 U3849 ( .A1(n3713), .A2(n2800), .B1(n402), .B2(n3281), .ZN(n2231)
         );
  OAI22_X1 U3850 ( .A1(n3713), .A2(n2813), .B1(n2812), .B2(n402), .ZN(n2244)
         );
  OAI22_X1 U3851 ( .A1(n3713), .A2(n2811), .B1(n2810), .B2(n402), .ZN(n2242)
         );
  OAI22_X1 U3852 ( .A1(n3713), .A2(n2831), .B1(n2830), .B2(n402), .ZN(n2262)
         );
  OAI22_X1 U3853 ( .A1(n3713), .A2(n2806), .B1(n2805), .B2(n402), .ZN(n2237)
         );
  OAI22_X1 U3854 ( .A1(n3713), .A2(n2807), .B1(n2806), .B2(n402), .ZN(n2238)
         );
  OAI22_X1 U3855 ( .A1(n3713), .A2(n2809), .B1(n2808), .B2(n402), .ZN(n2240)
         );
  OAI22_X1 U3856 ( .A1(n3713), .A2(n2810), .B1(n2809), .B2(n402), .ZN(n2241)
         );
  OAI22_X1 U3857 ( .A1(n3713), .A2(n2821), .B1(n2820), .B2(n402), .ZN(n2252)
         );
  OAI22_X1 U3858 ( .A1(n3713), .A2(n2822), .B1(n2821), .B2(n402), .ZN(n2253)
         );
  OAI22_X1 U3859 ( .A1(n3713), .A2(n2827), .B1(n2826), .B2(n402), .ZN(n2258)
         );
  OAI22_X1 U3860 ( .A1(n3713), .A2(n2823), .B1(n2822), .B2(n402), .ZN(n2254)
         );
  OAI22_X1 U3861 ( .A1(n3713), .A2(n2826), .B1(n2825), .B2(n402), .ZN(n2257)
         );
  OAI22_X1 U3862 ( .A1(n3713), .A2(n2818), .B1(n2817), .B2(n402), .ZN(n2249)
         );
  XNOR2_X1 U3863 ( .A(n1304), .B(n3656), .ZN(n1281) );
  XNOR2_X1 U3864 ( .A(n1283), .B(n1285), .ZN(n3656) );
  NAND2_X1 U3865 ( .A1(n1459), .A2(n1488), .ZN(n781) );
  OAI22_X1 U3866 ( .A1(n3667), .A2(n2983), .B1(n2982), .B2(n3571), .ZN(n2419)
         );
  OAI21_X1 U3867 ( .B1(n3680), .B2(n3738), .A(n3647), .ZN(n2400) );
  INV_X1 U3868 ( .A(n793), .ZN(n791) );
  NAND2_X1 U3869 ( .A1(n791), .A2(n794), .ZN(n561) );
  INV_X1 U3870 ( .A(n794), .ZN(n792) );
  NAND2_X2 U3871 ( .A1(n3747), .A2(n330), .ZN(n3660) );
  NAND2_X1 U3872 ( .A1(n3658), .A2(n3659), .ZN(n3661) );
  NAND2_X2 U3873 ( .A1(n3660), .A2(n3661), .ZN(n3746) );
  INV_X1 U3874 ( .A(n3747), .ZN(n3658) );
  INV_X4 U3875 ( .A(a[8]), .ZN(n3747) );
  OAI22_X1 U3876 ( .A1(n431), .A2(n3031), .B1(n381), .B2(n3288), .ZN(n2469) );
  BUF_X1 U3877 ( .A(n464), .Z(n3663) );
  INV_X8 U3878 ( .A(n3508), .ZN(n3664) );
  OAI21_X1 U3879 ( .B1(n3733), .B2(n3707), .A(n354), .ZN(n2230) );
  INV_X8 U3880 ( .A(n3705), .ZN(n408) );
  OAI21_X1 U3881 ( .B1(n3748), .B2(n3705), .A(n3574), .ZN(n2162) );
  NAND2_X1 U3882 ( .A1(n3460), .A2(n847), .ZN(n570) );
  OAI21_X1 U3883 ( .B1(n3753), .B2(n3746), .A(n3559), .ZN(n2468) );
  OAI21_X1 U3884 ( .B1(n3662), .B2(n3735), .A(n3731), .ZN(n2196) );
  OAI22_X1 U3885 ( .A1(n3670), .A2(n3158), .B1(n3157), .B2(n372), .ZN(n2599)
         );
  OAI22_X1 U3886 ( .A1(n3670), .A2(n3421), .B1(n3162), .B2(n372), .ZN(n2075)
         );
  OAI22_X1 U3887 ( .A1(n3670), .A2(n3159), .B1(n3158), .B2(n372), .ZN(n2600)
         );
  OAI22_X1 U3888 ( .A1(n3670), .A2(n3147), .B1(n3146), .B2(n372), .ZN(n2588)
         );
  OAI22_X1 U3889 ( .A1(n3670), .A2(n3160), .B1(n3159), .B2(n372), .ZN(n2601)
         );
  OAI22_X1 U3890 ( .A1(n3670), .A2(n3161), .B1(n3160), .B2(n372), .ZN(n2602)
         );
  OAI22_X1 U3891 ( .A1(n3670), .A2(n3157), .B1(n3156), .B2(n372), .ZN(n2598)
         );
  OAI22_X1 U3892 ( .A1(n3670), .A2(n3156), .B1(n3155), .B2(n372), .ZN(n2597)
         );
  OAI22_X1 U3893 ( .A1(n3670), .A2(n3155), .B1(n3154), .B2(n372), .ZN(n2596)
         );
  OAI22_X1 U3894 ( .A1(n3670), .A2(n3153), .B1(n3152), .B2(n372), .ZN(n2594)
         );
  OAI22_X1 U3895 ( .A1(n3670), .A2(n3152), .B1(n3151), .B2(n372), .ZN(n2593)
         );
  OAI22_X1 U3896 ( .A1(n3670), .A2(n3154), .B1(n3153), .B2(n372), .ZN(n2595)
         );
  OAI22_X1 U3897 ( .A1(n3670), .A2(n3142), .B1(n3141), .B2(n372), .ZN(n2583)
         );
  OAI22_X1 U3898 ( .A1(n3670), .A2(n3151), .B1(n3150), .B2(n372), .ZN(n2592)
         );
  OAI22_X1 U3899 ( .A1(n3670), .A2(n3148), .B1(n3147), .B2(n372), .ZN(n2589)
         );
  OAI22_X1 U3900 ( .A1(n3670), .A2(n3130), .B1(n372), .B2(n3421), .ZN(n2571)
         );
  OAI22_X1 U3901 ( .A1(n3670), .A2(n3138), .B1(n3137), .B2(n372), .ZN(n2579)
         );
  OAI22_X1 U3902 ( .A1(n3670), .A2(n3137), .B1(n3136), .B2(n372), .ZN(n2578)
         );
  OAI22_X1 U3903 ( .A1(n434), .A2(n3029), .B1(n3028), .B2(n3567), .ZN(n2466)
         );
  OAI22_X1 U3904 ( .A1(n3551), .A2(n3668), .B1(n3030), .B2(n3566), .ZN(n2071)
         );
  OAI22_X1 U3905 ( .A1(n3551), .A2(n3010), .B1(n3009), .B2(n3566), .ZN(n2447)
         );
  OAI22_X1 U3906 ( .A1(n3551), .A2(n3023), .B1(n3022), .B2(n3567), .ZN(n2460)
         );
  OAI22_X1 U3907 ( .A1(n3551), .A2(n3024), .B1(n3023), .B2(n3567), .ZN(n2461)
         );
  OAI22_X1 U3908 ( .A1(n3551), .A2(n3003), .B1(n3002), .B2(n3567), .ZN(n2440)
         );
  OAI22_X1 U3909 ( .A1(n3551), .A2(n3025), .B1(n3024), .B2(n3566), .ZN(n2462)
         );
  OAI22_X1 U3910 ( .A1(n3552), .A2(n3008), .B1(n3007), .B2(n3566), .ZN(n2445)
         );
  OAI22_X1 U3911 ( .A1(n3551), .A2(n3006), .B1(n3005), .B2(n3567), .ZN(n2443)
         );
  OAI22_X1 U3912 ( .A1(n434), .A2(n3017), .B1(n3016), .B2(n3566), .ZN(n2454)
         );
  OAI22_X1 U3913 ( .A1(n434), .A2(n3018), .B1(n3017), .B2(n3566), .ZN(n2455)
         );
  OAI22_X1 U3914 ( .A1(n3551), .A2(n3026), .B1(n3025), .B2(n3567), .ZN(n2463)
         );
  OAI22_X1 U3915 ( .A1(n434), .A2(n2998), .B1(n3567), .B2(n3668), .ZN(n2435)
         );
  BUF_X1 U3916 ( .A(n1283), .Z(n3666) );
  INV_X2 U3917 ( .A(n3668), .ZN(n3669) );
  OAI21_X1 U3918 ( .B1(n794), .B2(n788), .A(n789), .ZN(n787) );
  OAI21_X1 U3919 ( .B1(n3742), .B2(n3640), .A(n363), .ZN(n2128) );
  INV_X8 U3920 ( .A(n3671), .ZN(n3673) );
  INV_X8 U3921 ( .A(n3671), .ZN(n3672) );
  OAI21_X1 U3922 ( .B1(n531), .B2(n684), .A(n685), .ZN(n3674) );
  NAND2_X1 U3923 ( .A1(n3675), .A2(n3676), .ZN(n3678) );
  INV_X1 U3924 ( .A(n3749), .ZN(n3675) );
  INV_X1 U3925 ( .A(n324), .ZN(n3676) );
  OAI21_X1 U3926 ( .B1(n531), .B2(n684), .A(n685), .ZN(n683) );
  INV_X2 U3927 ( .A(n3686), .ZN(n685) );
  INV_X8 U3928 ( .A(n3696), .ZN(n396) );
  XNOR2_X1 U3929 ( .A(n595), .B(n3682), .ZN(product[63]) );
  XNOR2_X1 U3930 ( .A(n1042), .B(n1041), .ZN(n3682) );
  OAI22_X1 U3931 ( .A1(n3458), .A2(n2949), .B1(n2948), .B2(n3698), .ZN(n2384)
         );
  OAI21_X1 U3932 ( .B1(n3587), .B2(n3476), .A(n351), .ZN(n2264) );
  OAI21_X1 U3933 ( .B1(n3482), .B2(n3432), .A(n330), .ZN(n2502) );
  OAI21_X1 U3934 ( .B1(n3684), .B2(n3531), .A(n327), .ZN(n2536) );
  INV_X1 U3935 ( .A(n3456), .ZN(n1003) );
  INV_X4 U3936 ( .A(n3736), .ZN(n3683) );
  OAI22_X1 U3937 ( .A1(n3601), .A2(n3047), .B1(n3046), .B2(n381), .ZN(n2485)
         );
  INV_X1 U3938 ( .A(n431), .ZN(n3753) );
  AND2_X2 U3939 ( .A1(n3228), .A2(n3653), .ZN(n3685) );
  AOI21_X2 U3940 ( .B1(n706), .B2(n994), .A(n703), .ZN(n701) );
  OAI22_X1 U3941 ( .A1(n3712), .A2(n2808), .B1(n2807), .B2(n402), .ZN(n2239)
         );
  OAI22_X1 U3942 ( .A1(n3712), .A2(n2803), .B1(n2802), .B2(n402), .ZN(n2234)
         );
  OAI22_X1 U3943 ( .A1(n3712), .A2(n2801), .B1(n2800), .B2(n402), .ZN(n2232)
         );
  OAI22_X1 U3944 ( .A1(n3712), .A2(n2814), .B1(n2813), .B2(n402), .ZN(n2245)
         );
  OAI22_X1 U3945 ( .A1(n3712), .A2(n2802), .B1(n2801), .B2(n402), .ZN(n2233)
         );
  OAI22_X1 U3946 ( .A1(n3712), .A2(n3281), .B1(n2832), .B2(n402), .ZN(n2065)
         );
  OAI22_X1 U3947 ( .A1(n3712), .A2(n2824), .B1(n2823), .B2(n402), .ZN(n2255)
         );
  OAI22_X1 U3948 ( .A1(n3712), .A2(n2825), .B1(n2824), .B2(n402), .ZN(n2256)
         );
  OAI22_X1 U3949 ( .A1(n3712), .A2(n2820), .B1(n2819), .B2(n402), .ZN(n2251)
         );
  OAI22_X1 U3950 ( .A1(n3712), .A2(n2829), .B1(n2828), .B2(n402), .ZN(n2260)
         );
  OAI22_X1 U3951 ( .A1(n3712), .A2(n2828), .B1(n2827), .B2(n402), .ZN(n2259)
         );
  BUF_X1 U3952 ( .A(n687), .Z(n3686) );
  OAI21_X1 U3953 ( .B1(n3685), .B2(n3744), .A(n366), .ZN(n3754) );
  BUF_X1 U3954 ( .A(n612), .Z(n3687) );
  OAI21_X1 U3955 ( .B1(n3608), .B2(n707), .A(n708), .ZN(n3692) );
  AOI21_X2 U3956 ( .B1(n726), .B2(n709), .A(n710), .ZN(n708) );
  OAI22_X1 U3957 ( .A1(n428), .A2(n3067), .B1(n3066), .B2(n3664), .ZN(n2506)
         );
  INV_X1 U3958 ( .A(n3719), .ZN(n3694) );
  INV_X1 U3959 ( .A(n3694), .ZN(n3695) );
  NAND2_X1 U3960 ( .A1(n611), .A2(n981), .ZN(n604) );
  OAI22_X1 U3961 ( .A1(n446), .A2(n2877), .B1(n2876), .B2(n396), .ZN(n2310) );
  INV_X8 U3962 ( .A(n3697), .ZN(n3698) );
  INV_X1 U3963 ( .A(n3725), .ZN(n3699) );
  OAI21_X1 U3964 ( .B1(n3751), .B2(n3724), .A(n345), .ZN(n2332) );
  OAI21_X1 U3965 ( .B1(n3734), .B2(n3695), .A(n3669), .ZN(n2434) );
  OAI21_X1 U3966 ( .B1(n3736), .B2(n3696), .A(n348), .ZN(n2298) );
  OAI21_X1 U3967 ( .B1(n3743), .B2(n3700), .A(n342), .ZN(n2366) );
  OR2_X1 U3968 ( .A1(n1489), .A2(n1518), .ZN(n3701) );
  NOR2_X2 U3969 ( .A1(n788), .A2(n793), .ZN(n786) );
  NOR2_X2 U3970 ( .A1(n1489), .A2(n1518), .ZN(n788) );
  OAI21_X1 U3971 ( .B1(n807), .B2(n827), .A(n808), .ZN(n806) );
  XNOR2_X1 U3972 ( .A(n2572), .B(n3702), .ZN(n1571) );
  XNOR2_X1 U3973 ( .A(n2476), .B(n2540), .ZN(n3702) );
  BUF_X1 U3974 ( .A(n3487), .Z(n3703) );
  OAI21_X1 U3975 ( .B1(n3608), .B2(n604), .A(n605), .ZN(n603) );
  AOI21_X2 U3976 ( .B1(n761), .B2(n725), .A(n726), .ZN(n724) );
  INV_X2 U3977 ( .A(n3742), .ZN(n3720) );
  INV_X4 U3978 ( .A(n3681), .ZN(n372) );
  NAND2_X1 U3979 ( .A1(n1004), .A2(n778), .ZN(n558) );
  INV_X4 U3980 ( .A(n3707), .ZN(n402) );
  NAND2_X1 U3981 ( .A1(n1862), .A2(n1881), .ZN(n870) );
  OR2_X1 U3982 ( .A1(n1551), .A2(n1581), .ZN(n3708) );
  BUF_X1 U3983 ( .A(n3618), .Z(n3709) );
  INV_X1 U3984 ( .A(n798), .ZN(n796) );
  NAND2_X1 U3985 ( .A1(n798), .A2(n786), .ZN(n784) );
  OAI21_X1 U3986 ( .B1(n3608), .B2(n671), .A(n672), .ZN(n3711) );
  OAI21_X1 U3987 ( .B1(n531), .B2(n671), .A(n672), .ZN(n3710) );
  INV_X2 U3988 ( .A(n3733), .ZN(n3713) );
  INV_X1 U3989 ( .A(n3733), .ZN(n3712) );
  OAI21_X1 U3990 ( .B1(n531), .B2(n671), .A(n672), .ZN(n670) );
  INV_X1 U3991 ( .A(n3733), .ZN(n452) );
  NAND2_X1 U3992 ( .A1(n3666), .A2(n1304), .ZN(n3714) );
  NAND2_X1 U3993 ( .A1(n1304), .A2(n1285), .ZN(n3715) );
  NAND2_X1 U3994 ( .A1(n3666), .A2(n1285), .ZN(n3716) );
  NAND3_X1 U3995 ( .A1(n3714), .A2(n3716), .A3(n3715), .ZN(n1280) );
  NAND2_X1 U3996 ( .A1(n687), .A2(n673), .ZN(n3717) );
  INV_X1 U3997 ( .A(n676), .ZN(n3718) );
  AND2_X2 U3998 ( .A1(n3717), .A2(n3718), .ZN(n672) );
  NOR2_X1 U3999 ( .A1(n1259), .A2(n1280), .ZN(n735) );
  OAI21_X1 U4000 ( .B1(n677), .B2(n681), .A(n678), .ZN(n676) );
  XOR2_X1 U4001 ( .A(n805), .B(n563), .Z(product[32]) );
  OAI21_X1 U4002 ( .B1(n774), .B2(n3544), .A(n3473), .ZN(n771) );
  OAI21_X2 U4003 ( .B1(n805), .B2(n796), .A(n797), .ZN(n795) );
  OAI22_X1 U4004 ( .A1(n461), .A2(n2702), .B1(n2701), .B2(n3523), .ZN(n2130)
         );
  OAI22_X1 U4005 ( .A1(n461), .A2(n2705), .B1(n2704), .B2(n3523), .ZN(n2133)
         );
  OAI22_X1 U4006 ( .A1(n461), .A2(n2709), .B1(n2708), .B2(n3523), .ZN(n2137)
         );
  OAI22_X1 U4007 ( .A1(n461), .A2(n2708), .B1(n2707), .B2(n3523), .ZN(n2136)
         );
  OAI22_X1 U4008 ( .A1(n461), .A2(n2713), .B1(n2712), .B2(n3522), .ZN(n2141)
         );
  OAI22_X1 U4009 ( .A1(n461), .A2(n2721), .B1(n2720), .B2(n3523), .ZN(n2149)
         );
  OAI22_X1 U4010 ( .A1(n461), .A2(n2717), .B1(n2716), .B2(n3523), .ZN(n2145)
         );
  OAI22_X1 U4011 ( .A1(n461), .A2(n2719), .B1(n2718), .B2(n3523), .ZN(n2147)
         );
  OAI22_X1 U4012 ( .A1(n461), .A2(n2710), .B1(n2709), .B2(n3523), .ZN(n2138)
         );
  OAI22_X1 U4013 ( .A1(n461), .A2(n2725), .B1(n2724), .B2(n3522), .ZN(n2153)
         );
  OAI22_X1 U4014 ( .A1(n461), .A2(n2720), .B1(n2719), .B2(n3522), .ZN(n2148)
         );
  OAI22_X1 U4015 ( .A1(n461), .A2(n2724), .B1(n2723), .B2(n3522), .ZN(n2152)
         );
  OAI22_X1 U4016 ( .A1(n461), .A2(n2730), .B1(n2729), .B2(n3523), .ZN(n2158)
         );
  OAI22_X1 U4017 ( .A1(n3720), .A2(n2729), .B1(n2728), .B2(n3523), .ZN(n2157)
         );
  OAI22_X1 U4018 ( .A1(n3720), .A2(n2722), .B1(n2721), .B2(n3522), .ZN(n2150)
         );
  OAI22_X1 U4019 ( .A1(n3720), .A2(n2728), .B1(n2727), .B2(n3523), .ZN(n2156)
         );
  INV_X1 U4020 ( .A(n806), .ZN(n805) );
  NOR2_X2 U4021 ( .A1(n830), .A2(n842), .ZN(n828) );
  NAND2_X1 U4022 ( .A1(n1009), .A2(n804), .ZN(n563) );
  OAI21_X1 U4023 ( .B1(n805), .B2(n3575), .A(n804), .ZN(n802) );
  NOR2_X2 U4024 ( .A1(n772), .A2(n769), .ZN(n767) );
  NOR2_X2 U4025 ( .A1(n1403), .A2(n1430), .ZN(n772) );
  NAND2_X1 U4026 ( .A1(n809), .A2(n817), .ZN(n807) );
  INV_X1 U4027 ( .A(n3709), .ZN(n797) );
  INV_X1 U4028 ( .A(n3492), .ZN(n1010) );
  OAI21_X1 U4029 ( .B1(n815), .B2(n811), .A(n812), .ZN(n810) );
  NAND2_X1 U4030 ( .A1(n3445), .A2(n1641), .ZN(n812) );
  OAI22_X1 U4031 ( .A1(n422), .A2(n3133), .B1(n3132), .B2(n372), .ZN(n2574) );
  INV_X1 U4032 ( .A(n877), .ZN(n876) );
  INV_X1 U4033 ( .A(n3442), .ZN(n855) );
  AOI21_X2 U4034 ( .B1(n612), .B2(n981), .A(n607), .ZN(n605) );
  OAI22_X1 U4035 ( .A1(n452), .A2(n2815), .B1(n2814), .B2(n402), .ZN(n2246) );
  NAND2_X1 U4036 ( .A1(n1377), .A2(n1402), .ZN(n770) );
  NAND2_X1 U4037 ( .A1(n2572), .A2(n2476), .ZN(n3721) );
  NAND2_X1 U4038 ( .A1(n2572), .A2(n2540), .ZN(n3722) );
  NAND2_X1 U4039 ( .A1(n2476), .A2(n2540), .ZN(n3723) );
  NAND3_X1 U4040 ( .A1(n3721), .A2(n3723), .A3(n3722), .ZN(n1570) );
  OAI22_X1 U4041 ( .A1(n431), .A2(n3038), .B1(n3037), .B2(n381), .ZN(n2476) );
  OAI22_X1 U4042 ( .A1(n425), .A2(n3100), .B1(n3099), .B2(n3533), .ZN(n2540)
         );
  INV_X1 U4043 ( .A(n777), .ZN(n1004) );
  NOR2_X2 U4044 ( .A1(n780), .A2(n777), .ZN(n775) );
  OAI22_X1 U4045 ( .A1(n3595), .A2(n2752), .B1(n2751), .B2(n408), .ZN(n2181)
         );
  OAI22_X1 U4046 ( .A1(n3595), .A2(n2747), .B1(n2746), .B2(n408), .ZN(n2176)
         );
  OAI22_X1 U4047 ( .A1(n3595), .A2(n2741), .B1(n2740), .B2(n408), .ZN(n2170)
         );
  OAI22_X1 U4048 ( .A1(n3595), .A2(n2749), .B1(n2748), .B2(n408), .ZN(n2178)
         );
  OAI22_X1 U4049 ( .A1(n3595), .A2(n2745), .B1(n2744), .B2(n408), .ZN(n2174)
         );
  OAI22_X1 U4050 ( .A1(n3595), .A2(n2750), .B1(n2749), .B2(n408), .ZN(n2179)
         );
  OAI22_X1 U4051 ( .A1(n3595), .A2(n2746), .B1(n2745), .B2(n408), .ZN(n2175)
         );
  OAI22_X1 U4052 ( .A1(n3595), .A2(n2751), .B1(n2750), .B2(n408), .ZN(n2180)
         );
  OAI22_X1 U4053 ( .A1(n3595), .A2(n2748), .B1(n2747), .B2(n408), .ZN(n2177)
         );
  OAI22_X1 U4054 ( .A1(n3595), .A2(n2739), .B1(n2738), .B2(n408), .ZN(n2168)
         );
  OAI22_X1 U4055 ( .A1(n3595), .A2(n2755), .B1(n2754), .B2(n408), .ZN(n2184)
         );
  OAI22_X1 U4056 ( .A1(n3595), .A2(n2765), .B1(n2764), .B2(n408), .ZN(n2194)
         );
  OAI22_X1 U4057 ( .A1(n3595), .A2(n2757), .B1(n2756), .B2(n408), .ZN(n2186)
         );
  OAI22_X1 U4058 ( .A1(n3595), .A2(n3572), .B1(n2766), .B2(n408), .ZN(n2063)
         );
  OAI22_X1 U4059 ( .A1(n458), .A2(n2760), .B1(n2759), .B2(n408), .ZN(n2189) );
  OAI22_X1 U4060 ( .A1(n458), .A2(n2753), .B1(n2752), .B2(n408), .ZN(n2182) );
  OAI22_X1 U4061 ( .A1(n458), .A2(n2754), .B1(n2753), .B2(n408), .ZN(n2183) );
  OAI22_X1 U4062 ( .A1(n3595), .A2(n2756), .B1(n2755), .B2(n408), .ZN(n2185)
         );
  OAI22_X1 U4063 ( .A1(n458), .A2(n2761), .B1(n2760), .B2(n408), .ZN(n2190) );
  OAI22_X1 U4064 ( .A1(n458), .A2(n2762), .B1(n2761), .B2(n408), .ZN(n2191) );
  OAI22_X1 U4065 ( .A1(n458), .A2(n2759), .B1(n2758), .B2(n408), .ZN(n2188) );
  OAI22_X1 U4066 ( .A1(n458), .A2(n2764), .B1(n2763), .B2(n408), .ZN(n2193) );
  OAI22_X1 U4067 ( .A1(n458), .A2(n2758), .B1(n2757), .B2(n408), .ZN(n2187) );
  OAI22_X1 U4068 ( .A1(n458), .A2(n2763), .B1(n2762), .B2(n408), .ZN(n2192) );
  INV_X1 U4069 ( .A(n861), .ZN(n1018) );
  OAI21_X1 U4070 ( .B1(n861), .B2(n865), .A(n862), .ZN(n860) );
  NAND2_X1 U4071 ( .A1(n1820), .A2(n1841), .ZN(n862) );
  OAI21_X1 U4072 ( .B1(n3681), .B2(n3750), .A(n324), .ZN(n2570) );
  NAND2_X2 U4073 ( .A1(n1724), .A2(n1749), .ZN(n835) );
  AOI21_X2 U4074 ( .B1(n878), .B2(n897), .A(n879), .ZN(n877) );
  OAI21_X2 U4075 ( .B1(n898), .B2(n915), .A(n899), .ZN(n897) );
  NAND2_X1 U4076 ( .A1(n775), .A2(n767), .ZN(n765) );
  OAI22_X1 U4077 ( .A1(n3693), .A2(n3022), .B1(n3021), .B2(n3566), .ZN(n2459)
         );
  NOR2_X1 U4078 ( .A1(n1918), .A2(n1933), .ZN(n887) );
  NAND2_X2 U4079 ( .A1(n1918), .A2(n1933), .ZN(n888) );
  XOR2_X1 U4080 ( .A(n774), .B(n557), .Z(product[38]) );
  INV_X1 U4081 ( .A(n783), .ZN(n782) );
  AOI21_X1 U4082 ( .B1(n783), .B2(n3530), .A(n3419), .ZN(n774) );
  XNOR2_X1 U4083 ( .A(n650), .B(n539), .ZN(product[56]) );
  NAND2_X1 U4084 ( .A1(n1431), .A2(n1458), .ZN(n778) );
  XNOR2_X1 U4085 ( .A(n643), .B(n538), .ZN(product[57]) );
  OAI21_X1 U4086 ( .B1(n782), .B2(n3562), .A(n3629), .ZN(n779) );
  NAND2_X1 U4087 ( .A1(n1005), .A2(n3629), .ZN(n559) );
  OAI21_X1 U4088 ( .B1(n805), .B2(n784), .A(n3703), .ZN(n783) );
  OAI21_X1 U4089 ( .B1(n785), .B2(n765), .A(n766), .ZN(n764) );
  INV_X1 U4090 ( .A(n3612), .ZN(n826) );
  AOI21_X2 U4091 ( .B1(n683), .B2(n631), .A(n632), .ZN(n630) );
  XNOR2_X1 U4092 ( .A(n717), .B(n549), .ZN(product[46]) );
  XNOR2_X1 U4093 ( .A(n662), .B(n541), .ZN(product[54]) );
  INV_X1 U4094 ( .A(n3429), .ZN(n726) );
  OAI21_X1 U4095 ( .B1(n3429), .B2(n613), .A(n614), .ZN(n612) );
  OAI21_X1 U4096 ( .B1(n731), .B2(n748), .A(n732), .ZN(n730) );
  XNOR2_X1 U4097 ( .A(n698), .B(n546), .ZN(product[49]) );
  XNOR2_X1 U4098 ( .A(n737), .B(n551), .ZN(product[44]) );
  XNOR2_X1 U4099 ( .A(n623), .B(n536), .ZN(product[59]) );
  NAND2_X1 U4100 ( .A1(n763), .A2(n806), .ZN(n3727) );
  INV_X1 U4101 ( .A(n764), .ZN(n3728) );
  INV_X1 U4102 ( .A(n3748), .ZN(n3729) );
  INV_X2 U4103 ( .A(n3730), .ZN(n3731) );
  AOI21_X1 U4104 ( .B1(n3641), .B2(n654), .A(n655), .ZN(n653) );
  NOR2_X1 U4105 ( .A1(n784), .A2(n765), .ZN(n763) );
  XOR2_X1 U4106 ( .A(n724), .B(n550), .Z(product[45]) );
  OAI21_X1 U4107 ( .B1(n724), .B2(n718), .A(n719), .ZN(n717) );
  AOI21_X1 U4108 ( .B1(n3704), .B2(n980), .A(n600), .ZN(n3732) );
  OAI22_X1 U4109 ( .A1(n3623), .A2(n2914), .B1(n2913), .B2(n393), .ZN(n2348)
         );
  AND2_X2 U4110 ( .A1(n3232), .A2(n3545), .ZN(n3733) );
  INV_X4 U4111 ( .A(n3734), .ZN(n434) );
  AND2_X2 U4112 ( .A1(n3234), .A2(n3550), .ZN(n3736) );
  OAI22_X1 U4113 ( .A1(n446), .A2(n2883), .B1(n2882), .B2(n396), .ZN(n2316) );
  OAI22_X1 U4114 ( .A1(n455), .A2(n2789), .B1(n2788), .B2(n3630), .ZN(n2219)
         );
  XNOR2_X2 U4115 ( .A(n3741), .B(n348), .ZN(n3740) );
  INV_X4 U4116 ( .A(n3742), .ZN(n461) );
  INV_X8 U4117 ( .A(n3746), .ZN(n381) );
  INV_X4 U4118 ( .A(n3748), .ZN(n458) );
  INV_X4 U4119 ( .A(n3750), .ZN(n422) );
  AOI21_X2 U4120 ( .B1(n670), .B2(n989), .A(n667), .ZN(n665) );
  XOR2_X1 U4121 ( .A(n665), .B(n542), .Z(product[53]) );
  OAI21_X1 U4122 ( .B1(n665), .B2(n663), .A(n664), .ZN(n662) );
  OAI21_X1 U4123 ( .B1(n630), .B2(n624), .A(n625), .ZN(n623) );
  XOR2_X1 U4124 ( .A(n630), .B(n537), .Z(product[58]) );
  XNOR2_X1 U4125 ( .A(n3603), .B(n553), .ZN(product[42]) );
  OAI21_X1 U4126 ( .B1(n744), .B2(n738), .A(n739), .ZN(n737) );
  XOR2_X1 U4127 ( .A(n3560), .B(n552), .Z(product[43]) );
  XNOR2_X1 U4128 ( .A(n3692), .B(n548), .ZN(product[47]) );
  OAI21_X1 U4129 ( .B1(n701), .B2(n699), .A(n700), .ZN(n698) );
  XOR2_X1 U4130 ( .A(n701), .B(n547), .Z(product[48]) );
  OAI22_X1 U4131 ( .A1(n3670), .A2(n3131), .B1(n3130), .B2(n372), .ZN(n2572)
         );
  XNOR2_X1 U4132 ( .A(n3600), .B(n555), .ZN(product[40]) );
  AOI21_X1 U4133 ( .B1(n3557), .B2(n757), .A(n758), .ZN(n756) );
  AOI21_X1 U4134 ( .B1(n3557), .B2(n611), .A(n3687), .ZN(n610) );
  INV_X4 U4135 ( .A(n3751), .ZN(n443) );
  XNOR2_X1 U4136 ( .A(n3704), .B(n534), .ZN(product[61]) );
  XNOR2_X1 U4137 ( .A(n3711), .B(n543), .ZN(product[52]) );
  OAI21_X1 U4138 ( .B1(n3726), .B2(n651), .A(n652), .ZN(n650) );
  OAI21_X1 U4139 ( .B1(n653), .B2(n644), .A(n645), .ZN(n643) );
  XOR2_X1 U4140 ( .A(n3726), .B(n540), .Z(product[55]) );
  INV_X1 U4141 ( .A(n3608), .ZN(n761) );
  OAI21_X1 U4142 ( .B1(n531), .B2(n707), .A(n708), .ZN(n706) );
  OAI21_X1 U4143 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  INV_X2 U4144 ( .A(n594), .ZN(product[1]) );
  INV_X2 U4145 ( .A(n699), .ZN(n993) );
  INV_X2 U4146 ( .A(n680), .ZN(n991) );
  INV_X2 U4147 ( .A(n677), .ZN(n990) );
  INV_X2 U4148 ( .A(n663), .ZN(n988) );
  INV_X2 U4149 ( .A(n660), .ZN(n987) );
  INV_X2 U4150 ( .A(n651), .ZN(n986) );
  INV_X2 U4151 ( .A(n648), .ZN(n985) );
  INV_X2 U4152 ( .A(n596), .ZN(n979) );
  INV_X2 U4153 ( .A(n978), .ZN(n976) );
  INV_X2 U4154 ( .A(n975), .ZN(n973) );
  INV_X2 U4155 ( .A(n967), .ZN(n965) );
  INV_X2 U4156 ( .A(n959), .ZN(n957) );
  INV_X2 U4157 ( .A(n955), .ZN(n954) );
  INV_X2 U4158 ( .A(n953), .ZN(n951) );
  INV_X2 U4159 ( .A(n948), .ZN(n946) );
  INV_X2 U4160 ( .A(n941), .ZN(n939) );
  INV_X2 U4161 ( .A(n937), .ZN(n936) );
  INV_X2 U4162 ( .A(n935), .ZN(n933) );
  INV_X2 U4163 ( .A(n930), .ZN(n928) );
  INV_X2 U4164 ( .A(n924), .ZN(n923) );
  INV_X2 U4165 ( .A(n915), .ZN(n914) );
  INV_X2 U4166 ( .A(n913), .ZN(n911) );
  INV_X2 U4167 ( .A(n903), .ZN(n901) );
  INV_X2 U4168 ( .A(n891), .ZN(n893) );
  INV_X2 U4169 ( .A(n888), .ZN(n886) );
  INV_X2 U4170 ( .A(n875), .ZN(n873) );
  INV_X2 U4171 ( .A(n835), .ZN(n833) );
  INV_X2 U4172 ( .A(n825), .ZN(n823) );
  INV_X2 U4173 ( .A(n752), .ZN(n750) );
  INV_X2 U4174 ( .A(n748), .ZN(n746) );
  INV_X2 U4175 ( .A(n736), .ZN(n734) );
  INV_X2 U4176 ( .A(n719), .ZN(n721) );
  INV_X2 U4177 ( .A(n718), .ZN(n996) );
  INV_X2 U4178 ( .A(n716), .ZN(n714) );
  INV_X2 U4179 ( .A(n715), .ZN(n995) );
  INV_X2 U4180 ( .A(n712), .ZN(n710) );
  INV_X2 U4181 ( .A(n711), .ZN(n709) );
  INV_X2 U4182 ( .A(n705), .ZN(n703) );
  INV_X2 U4183 ( .A(n704), .ZN(n994) );
  INV_X2 U4184 ( .A(n691), .ZN(n689) );
  INV_X2 U4185 ( .A(n686), .ZN(n684) );
  INV_X2 U4186 ( .A(n3674), .ZN(n682) );
  INV_X2 U4187 ( .A(n669), .ZN(n667) );
  INV_X2 U4188 ( .A(n668), .ZN(n989) );
  INV_X2 U4189 ( .A(n656), .ZN(n654) );
  INV_X2 U4190 ( .A(n647), .ZN(n645) );
  INV_X2 U4191 ( .A(n646), .ZN(n644) );
  INV_X2 U4192 ( .A(n642), .ZN(n640) );
  INV_X2 U4193 ( .A(n641), .ZN(n984) );
  INV_X2 U4194 ( .A(n634), .ZN(n632) );
  INV_X2 U4195 ( .A(n633), .ZN(n631) );
  INV_X2 U4196 ( .A(n625), .ZN(n627) );
  INV_X2 U4197 ( .A(n624), .ZN(n983) );
  INV_X2 U4198 ( .A(n622), .ZN(n620) );
  INV_X2 U4199 ( .A(n621), .ZN(n982) );
  INV_X2 U4200 ( .A(n609), .ZN(n607) );
  INV_X2 U4201 ( .A(n608), .ZN(n981) );
  INV_X2 U4202 ( .A(n602), .ZN(n600) );
  INV_X2 U4203 ( .A(n601), .ZN(n980) );
  INV_X2 U4204 ( .A(n3559), .ZN(n3288) );
  INV_X2 U4205 ( .A(n3647), .ZN(n3286) );
  INV_X2 U4206 ( .A(n348), .ZN(n3283) );
  INV_X2 U4207 ( .A(n351), .ZN(n3282) );
  NAND2_X2 U4208 ( .A1(n321), .A2(n3752), .ZN(n3195) );
  NAND2_X2 U4209 ( .A1(n324), .A2(n3752), .ZN(n3162) );
  NAND2_X2 U4210 ( .A1(n327), .A2(n3752), .ZN(n3129) );
  NAND2_X2 U4211 ( .A1(n330), .A2(n3752), .ZN(n3096) );
  NAND2_X2 U4212 ( .A1(n3559), .A2(n3752), .ZN(n3063) );
  NAND2_X2 U4213 ( .A1(n3669), .A2(n3752), .ZN(n3030) );
  NAND2_X2 U4214 ( .A1(n3647), .A2(n3752), .ZN(n2997) );
  NAND2_X2 U4215 ( .A1(n342), .A2(n3752), .ZN(n2964) );
  NAND2_X2 U4216 ( .A1(n345), .A2(n3752), .ZN(n2931) );
  NAND2_X2 U4217 ( .A1(n348), .A2(n3752), .ZN(n2898) );
  NAND2_X2 U4218 ( .A1(n351), .A2(n3752), .ZN(n2865) );
  NAND2_X2 U4219 ( .A1(n354), .A2(n3752), .ZN(n2832) );
  NAND2_X2 U4220 ( .A1(n3731), .A2(n3752), .ZN(n2799) );
  NAND2_X2 U4221 ( .A1(n3574), .A2(n3752), .ZN(n2766) );
  NAND2_X2 U4222 ( .A1(n363), .A2(n3752), .ZN(n2733) );
  NAND2_X2 U4223 ( .A1(n366), .A2(n3752), .ZN(n2700) );
  NOR2_X2 U4224 ( .A1(n372), .A2(n3752), .ZN(n2603) );
  NOR2_X2 U4225 ( .A1(n3533), .A2(n3752), .ZN(n2569) );
  NOR2_X2 U4226 ( .A1(n3664), .A2(n3752), .ZN(n2535) );
  NOR2_X2 U4227 ( .A1(n381), .A2(n3752), .ZN(n2501) );
  NOR2_X2 U4228 ( .A1(n3566), .A2(n3752), .ZN(n2467) );
  NOR2_X2 U4229 ( .A1(n3571), .A2(n3752), .ZN(n2433) );
  NOR2_X2 U4230 ( .A1(n3698), .A2(n3752), .ZN(n2399) );
  NOR2_X2 U4231 ( .A1(n393), .A2(n3752), .ZN(n2365) );
  NOR2_X2 U4232 ( .A1(n396), .A2(n3752), .ZN(n2331) );
  NOR2_X2 U4233 ( .A1(n3673), .A2(n3752), .ZN(n2297) );
  NOR2_X2 U4234 ( .A1(n402), .A2(n3752), .ZN(n2263) );
  NOR2_X2 U4235 ( .A1(n3630), .A2(n3752), .ZN(n2229) );
  NOR2_X2 U4236 ( .A1(n408), .A2(n3752), .ZN(n2195) );
  NOR2_X2 U4237 ( .A1(n3522), .A2(n3752), .ZN(n2161) );
  NOR2_X2 U4238 ( .A1(n3655), .A2(n3752), .ZN(n2127) );
  INV_X2 U4239 ( .A(n1548), .ZN(n1580) );
  INV_X2 U4240 ( .A(n1374), .ZN(n1375) );
  INV_X2 U4241 ( .A(n1324), .ZN(n1325) );
  INV_X2 U4242 ( .A(n1278), .ZN(n1279) );
  INV_X2 U4243 ( .A(n1236), .ZN(n1237) );
  INV_X2 U4244 ( .A(n1198), .ZN(n1199) );
  INV_X2 U4245 ( .A(n1164), .ZN(n1165) );
  INV_X2 U4246 ( .A(n1134), .ZN(n1135) );
  INV_X2 U4247 ( .A(n1108), .ZN(n1109) );
  INV_X2 U4248 ( .A(n1086), .ZN(n1087) );
  INV_X2 U4249 ( .A(n1068), .ZN(n1069) );
  INV_X2 U4250 ( .A(n1054), .ZN(n1055) );
  INV_X2 U4251 ( .A(n1044), .ZN(n1045) );
  XOR2_X1 U4252 ( .A(n3754), .B(n3755), .Z(n1041) );
  XOR2_X1 U4253 ( .A(n2077), .B(n1044), .Z(n3755) );
  INV_X2 U4254 ( .A(n977), .ZN(n1040) );
  INV_X2 U4255 ( .A(n974), .ZN(n972) );
  INV_X2 U4256 ( .A(n969), .ZN(n1038) );
  INV_X2 U4257 ( .A(n966), .ZN(n964) );
  INV_X2 U4258 ( .A(n961), .ZN(n1036) );
  INV_X2 U4259 ( .A(n958), .ZN(n956) );
  INV_X2 U4260 ( .A(n952), .ZN(n950) );
  INV_X2 U4261 ( .A(n947), .ZN(n945) );
  INV_X2 U4262 ( .A(n940), .ZN(n938) );
  INV_X2 U4263 ( .A(n934), .ZN(n932) );
  INV_X2 U4264 ( .A(n929), .ZN(n927) );
  INV_X2 U4265 ( .A(n921), .ZN(n1029) );
  INV_X2 U4266 ( .A(n918), .ZN(n1028) );
  INV_X2 U4267 ( .A(n912), .ZN(n910) );
  INV_X2 U4268 ( .A(n902), .ZN(n900) );
  INV_X2 U4269 ( .A(n890), .ZN(n892) );
  INV_X2 U4270 ( .A(n880), .ZN(n1022) );
  INV_X2 U4271 ( .A(n874), .ZN(n872) );
  INV_X2 U4272 ( .A(n869), .ZN(n1020) );
  INV_X2 U4273 ( .A(n849), .ZN(n851) );
  INV_X2 U4274 ( .A(n759), .ZN(n757) );
endmodule


module mul32_2_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n321, n324, n327, n330, n333, n336, n339, n342, n345, n348, n351,
         n354, n357, n360, n363, n366, n369, n372, n375, n378, n381, n384,
         n387, n390, n396, n399, n402, n405, n408, n411, n414, n416, n419,
         n422, n428, n434, n437, n440, n443, n446, n449, n452, n455, n458,
         n461, n464, n465, n469, n471, n473, n475, n477, n479, n481, n483,
         n485, n487, n489, n491, n493, n495, n497, n499, n501, n503, n505,
         n507, n509, n511, n513, n515, n517, n519, n521, n523, n525, n527,
         n529, n531, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n600, n601, n602, n603, n604, n605, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n620, n621, n622,
         n623, n624, n625, n627, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n667, n668, n669, n670, n671,
         n672, n673, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n714, n715, n716, n717, n718, n719,
         n721, n724, n726, n727, n728, n729, n730, n731, n732, n734, n735,
         n736, n737, n738, n739, n741, n744, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n763, n764, n765, n766, n768, n769, n770, n771, n772, n773, n774,
         n775, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n838, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n999, n1000, n1003, n1005,
         n1006, n1008, n1009, n1010, n1011, n1012, n1018, n1019, n1020, n1022,
         n1026, n1028, n1029, n1036, n1038, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3240, n3242, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3290, n3292, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761;
  assign n321 = a[1];
  assign n324 = a[3];
  assign n327 = a[5];
  assign n330 = a[7];
  assign n333 = a[9];
  assign n336 = a[11];
  assign n339 = a[13];
  assign n342 = a[15];
  assign n345 = a[17];
  assign n348 = a[19];
  assign n351 = a[21];
  assign n354 = a[23];
  assign n357 = a[25];
  assign n360 = a[27];
  assign n363 = a[29];
  assign n366 = a[31];
  assign n465 = b[0];
  assign n469 = b[1];
  assign n471 = b[2];
  assign n473 = b[3];
  assign n475 = b[4];
  assign n477 = b[5];
  assign n479 = b[6];
  assign n481 = b[7];
  assign n483 = b[8];
  assign n485 = b[9];
  assign n487 = b[10];
  assign n489 = b[11];
  assign n491 = b[12];
  assign n493 = b[13];
  assign n495 = b[14];
  assign n497 = b[15];
  assign n499 = b[16];
  assign n501 = b[17];
  assign n503 = b[18];
  assign n505 = b[19];
  assign n507 = b[20];
  assign n509 = b[21];
  assign n511 = b[22];
  assign n513 = b[23];
  assign n515 = b[24];
  assign n517 = b[25];
  assign n519 = b[26];
  assign n521 = b[27];
  assign n523 = b[28];
  assign n525 = b[29];
  assign n527 = b[30];
  assign n529 = b[31];

  NAND2_X4 U322 ( .A1(n979), .A2(n597), .ZN(n533) );
  NOR2_X4 U324 ( .A1(n1043), .A2(n1046), .ZN(n596) );
  NAND2_X4 U325 ( .A1(n1043), .A2(n1046), .ZN(n597) );
  NAND2_X4 U330 ( .A1(n980), .A2(n602), .ZN(n534) );
  NOR2_X4 U332 ( .A1(n1050), .A2(n1047), .ZN(n601) );
  NAND2_X4 U333 ( .A1(n1050), .A2(n1047), .ZN(n602) );
  XOR2_X2 U334 ( .A(n610), .B(n535), .Z(product[60]) );
  NAND2_X4 U340 ( .A1(n981), .A2(n609), .ZN(n535) );
  NOR2_X4 U342 ( .A1(n1051), .A2(n1056), .ZN(n608) );
  NAND2_X4 U343 ( .A1(n1051), .A2(n1056), .ZN(n609) );
  NOR2_X4 U350 ( .A1(n633), .A2(n617), .ZN(n615) );
  NAND2_X4 U352 ( .A1(n983), .A2(n982), .ZN(n617) );
  AOI21_X4 U353 ( .B1(n982), .B2(n627), .A(n620), .ZN(n618) );
  NAND2_X4 U356 ( .A1(n982), .A2(n622), .ZN(n536) );
  NOR2_X4 U358 ( .A1(n1057), .A2(n1062), .ZN(n621) );
  NAND2_X4 U359 ( .A1(n1057), .A2(n1062), .ZN(n622) );
  NAND2_X4 U366 ( .A1(n983), .A2(n625), .ZN(n537) );
  NOR2_X4 U368 ( .A1(n1063), .A2(n1070), .ZN(n624) );
  NAND2_X4 U369 ( .A1(n1063), .A2(n1070), .ZN(n625) );
  NAND2_X4 U374 ( .A1(n673), .A2(n635), .ZN(n633) );
  NOR2_X4 U376 ( .A1(n656), .A2(n637), .ZN(n635) );
  OAI21_X4 U377 ( .B1(n657), .B2(n637), .A(n638), .ZN(n636) );
  NAND2_X4 U378 ( .A1(n646), .A2(n984), .ZN(n637) );
  AOI21_X4 U379 ( .B1(n647), .B2(n984), .A(n640), .ZN(n638) );
  NAND2_X4 U382 ( .A1(n984), .A2(n642), .ZN(n538) );
  NOR2_X4 U384 ( .A1(n1071), .A2(n1078), .ZN(n641) );
  NAND2_X4 U385 ( .A1(n1071), .A2(n1078), .ZN(n642) );
  NOR2_X4 U390 ( .A1(n651), .A2(n648), .ZN(n646) );
  OAI21_X4 U391 ( .B1(n648), .B2(n652), .A(n649), .ZN(n647) );
  NAND2_X4 U392 ( .A1(n985), .A2(n649), .ZN(n539) );
  NOR2_X4 U394 ( .A1(n1079), .A2(n1088), .ZN(n648) );
  NAND2_X4 U395 ( .A1(n1079), .A2(n1088), .ZN(n649) );
  NAND2_X4 U398 ( .A1(n986), .A2(n652), .ZN(n540) );
  NOR2_X4 U400 ( .A1(n1089), .A2(n1098), .ZN(n651) );
  NAND2_X4 U401 ( .A1(n1089), .A2(n1098), .ZN(n652) );
  NAND2_X4 U406 ( .A1(n658), .A2(n989), .ZN(n656) );
  AOI21_X4 U407 ( .B1(n658), .B2(n667), .A(n659), .ZN(n657) );
  NOR2_X4 U408 ( .A1(n663), .A2(n660), .ZN(n658) );
  OAI21_X4 U409 ( .B1(n660), .B2(n664), .A(n661), .ZN(n659) );
  NAND2_X4 U410 ( .A1(n987), .A2(n661), .ZN(n541) );
  NOR2_X4 U412 ( .A1(n1099), .A2(n1110), .ZN(n660) );
  NAND2_X4 U413 ( .A1(n1099), .A2(n1110), .ZN(n661) );
  NAND2_X4 U416 ( .A1(n988), .A2(n664), .ZN(n542) );
  NOR2_X4 U418 ( .A1(n1111), .A2(n1122), .ZN(n663) );
  NAND2_X4 U419 ( .A1(n1111), .A2(n1122), .ZN(n664) );
  NAND2_X4 U424 ( .A1(n989), .A2(n669), .ZN(n543) );
  XNOR2_X2 U428 ( .A(n679), .B(n544), .ZN(product[51]) );
  NOR2_X4 U434 ( .A1(n680), .A2(n677), .ZN(n673) );
  OAI21_X4 U435 ( .B1(n677), .B2(n681), .A(n678), .ZN(n676) );
  NAND2_X4 U436 ( .A1(n990), .A2(n678), .ZN(n544) );
  NOR2_X4 U438 ( .A1(n1137), .A2(n1150), .ZN(n677) );
  NAND2_X4 U439 ( .A1(n1137), .A2(n1150), .ZN(n678) );
  NAND2_X4 U442 ( .A1(n991), .A2(n681), .ZN(n545) );
  NOR2_X4 U444 ( .A1(n1151), .A2(n1166), .ZN(n680) );
  NAND2_X4 U445 ( .A1(n1151), .A2(n1166), .ZN(n681) );
  NOR2_X4 U455 ( .A1(n692), .A2(n711), .ZN(n690) );
  OAI21_X4 U456 ( .B1(n692), .B2(n712), .A(n693), .ZN(n691) );
  OAI21_X4 U460 ( .B1(n696), .B2(n700), .A(n697), .ZN(n695) );
  NAND2_X4 U461 ( .A1(n992), .A2(n697), .ZN(n546) );
  NOR2_X4 U463 ( .A1(n1167), .A2(n1182), .ZN(n696) );
  NAND2_X4 U464 ( .A1(n1167), .A2(n1182), .ZN(n697) );
  NOR2_X4 U469 ( .A1(n1183), .A2(n1200), .ZN(n699) );
  NAND2_X4 U470 ( .A1(n1183), .A2(n1200), .ZN(n700) );
  NAND2_X4 U475 ( .A1(n994), .A2(n705), .ZN(n548) );
  NOR2_X4 U477 ( .A1(n1201), .A2(n1218), .ZN(n704) );
  NAND2_X4 U478 ( .A1(n1201), .A2(n1218), .ZN(n705) );
  NAND2_X4 U481 ( .A1(n3485), .A2(n709), .ZN(n707) );
  NAND2_X4 U499 ( .A1(n996), .A2(n719), .ZN(n550) );
  NOR2_X4 U501 ( .A1(n1239), .A2(n1258), .ZN(n718) );
  NAND2_X4 U502 ( .A1(n1239), .A2(n1258), .ZN(n719) );
  NAND2_X4 U525 ( .A1(n3655), .A2(n739), .ZN(n552) );
  NAND2_X4 U533 ( .A1(n999), .A2(n748), .ZN(n553) );
  XOR2_X2 U537 ( .A(n756), .B(n554), .Z(product[41]) );
  NAND2_X4 U543 ( .A1(n1000), .A2(n755), .ZN(n554) );
  XNOR2_X2 U574 ( .A(n779), .B(n558), .ZN(product[37]) );
  XOR2_X2 U582 ( .A(n782), .B(n559), .Z(product[36]) );
  XOR2_X2 U588 ( .A(n790), .B(n560), .Z(product[35]) );
  XNOR2_X2 U607 ( .A(n802), .B(n562), .ZN(product[33]) );
  NOR2_X4 U615 ( .A1(n1551), .A2(n1581), .ZN(n800) );
  XNOR2_X2 U623 ( .A(n813), .B(n564), .ZN(product[31]) );
  NAND2_X4 U630 ( .A1(n1010), .A2(n812), .ZN(n564) );
  XOR2_X2 U634 ( .A(n816), .B(n565), .Z(product[30]) );
  XOR2_X2 U640 ( .A(n821), .B(n566), .Z(product[29]) );
  XNOR2_X2 U648 ( .A(n826), .B(n567), .ZN(product[28]) );
  AOI21_X4 U649 ( .B1(n826), .B2(n822), .A(n823), .ZN(n821) );
  XOR2_X2 U656 ( .A(n836), .B(n568), .Z(product[27]) );
  XNOR2_X2 U669 ( .A(n841), .B(n569), .ZN(product[26]) );
  AOI21_X4 U670 ( .B1(n841), .B2(n3480), .A(n838), .ZN(n836) );
  XNOR2_X2 U677 ( .A(n848), .B(n570), .ZN(product[25]) );
  XOR2_X2 U687 ( .A(n855), .B(n571), .Z(product[24]) );
  XNOR2_X2 U697 ( .A(n863), .B(n572), .ZN(product[23]) );
  NAND2_X4 U704 ( .A1(n1018), .A2(n862), .ZN(n572) );
  XOR2_X2 U708 ( .A(n866), .B(n573), .Z(product[22]) );
  OAI21_X4 U709 ( .B1(n866), .B2(n864), .A(n865), .ZN(n863) );
  NAND2_X4 U710 ( .A1(n1019), .A2(n865), .ZN(n573) );
  NOR2_X4 U712 ( .A1(n1842), .A2(n1861), .ZN(n864) );
  XOR2_X2 U714 ( .A(n871), .B(n574), .Z(product[21]) );
  AOI21_X4 U715 ( .B1(n876), .B2(n867), .A(n868), .ZN(n866) );
  NOR2_X4 U716 ( .A1(n869), .A2(n874), .ZN(n867) );
  OAI21_X4 U717 ( .B1(n869), .B2(n875), .A(n870), .ZN(n868) );
  NAND2_X4 U718 ( .A1(n1020), .A2(n870), .ZN(n574) );
  NOR2_X4 U720 ( .A1(n1862), .A2(n1881), .ZN(n869) );
  XNOR2_X2 U722 ( .A(n876), .B(n575), .ZN(product[20]) );
  AOI21_X4 U723 ( .B1(n876), .B2(n872), .A(n873), .ZN(n871) );
  NAND2_X4 U726 ( .A1(n872), .A2(n875), .ZN(n575) );
  XNOR2_X2 U730 ( .A(n882), .B(n576), .ZN(product[19]) );
  NOR2_X4 U733 ( .A1(n883), .A2(n880), .ZN(n878) );
  NAND2_X4 U735 ( .A1(n1022), .A2(n881), .ZN(n576) );
  NOR2_X4 U737 ( .A1(n1900), .A2(n1917), .ZN(n880) );
  XNOR2_X2 U739 ( .A(n889), .B(n577), .ZN(product[18]) );
  NAND2_X4 U741 ( .A1(n885), .A2(n892), .ZN(n883) );
  NAND2_X4 U745 ( .A1(n885), .A2(n888), .ZN(n577) );
  XOR2_X2 U749 ( .A(n896), .B(n578), .Z(product[17]) );
  OAI21_X4 U750 ( .B1(n896), .B2(n890), .A(n891), .ZN(n889) );
  NAND2_X4 U755 ( .A1(n892), .A2(n891), .ZN(n578) );
  NOR2_X4 U757 ( .A1(n1934), .A2(n1949), .ZN(n890) );
  NAND2_X4 U758 ( .A1(n1934), .A2(n1949), .ZN(n891) );
  XOR2_X2 U759 ( .A(n904), .B(n579), .Z(product[16]) );
  OAI21_X4 U761 ( .B1(n898), .B2(n915), .A(n899), .ZN(n897) );
  NAND2_X4 U762 ( .A1(n905), .A2(n900), .ZN(n898) );
  NAND2_X4 U766 ( .A1(n900), .A2(n903), .ZN(n579) );
  NOR2_X4 U768 ( .A1(n1950), .A2(n1963), .ZN(n902) );
  NAND2_X4 U769 ( .A1(n1950), .A2(n1963), .ZN(n903) );
  XOR2_X2 U770 ( .A(n909), .B(n580), .Z(product[15]) );
  NOR2_X4 U772 ( .A1(n907), .A2(n912), .ZN(n905) );
  NAND2_X4 U774 ( .A1(n1026), .A2(n908), .ZN(n580) );
  NOR2_X4 U776 ( .A1(n1964), .A2(n1977), .ZN(n907) );
  XNOR2_X2 U778 ( .A(n914), .B(n581), .ZN(product[14]) );
  AOI21_X4 U779 ( .B1(n914), .B2(n910), .A(n911), .ZN(n909) );
  NAND2_X4 U782 ( .A1(n910), .A2(n913), .ZN(n581) );
  NOR2_X4 U784 ( .A1(n1978), .A2(n1989), .ZN(n912) );
  NAND2_X4 U785 ( .A1(n1978), .A2(n1989), .ZN(n913) );
  XNOR2_X2 U786 ( .A(n920), .B(n582), .ZN(product[13]) );
  AOI21_X4 U788 ( .B1(n916), .B2(n924), .A(n917), .ZN(n915) );
  NOR2_X4 U789 ( .A1(n918), .A2(n921), .ZN(n916) );
  OAI21_X4 U790 ( .B1(n918), .B2(n922), .A(n919), .ZN(n917) );
  NAND2_X4 U791 ( .A1(n1028), .A2(n919), .ZN(n582) );
  NOR2_X4 U793 ( .A1(n1990), .A2(n2001), .ZN(n918) );
  NAND2_X4 U794 ( .A1(n1990), .A2(n2001), .ZN(n919) );
  XOR2_X2 U795 ( .A(n923), .B(n583), .Z(product[12]) );
  OAI21_X4 U796 ( .B1(n923), .B2(n921), .A(n922), .ZN(n920) );
  NAND2_X4 U797 ( .A1(n1029), .A2(n922), .ZN(n583) );
  NOR2_X4 U799 ( .A1(n2002), .A2(n2011), .ZN(n921) );
  NAND2_X4 U800 ( .A1(n2002), .A2(n2011), .ZN(n922) );
  XOR2_X2 U801 ( .A(n931), .B(n584), .Z(product[11]) );
  OAI21_X4 U803 ( .B1(n925), .B2(n937), .A(n926), .ZN(n924) );
  NAND2_X4 U804 ( .A1(n932), .A2(n927), .ZN(n925) );
  AOI21_X4 U805 ( .B1(n927), .B2(n933), .A(n928), .ZN(n926) );
  NAND2_X4 U808 ( .A1(n927), .A2(n930), .ZN(n584) );
  NOR2_X4 U810 ( .A1(n2012), .A2(n2021), .ZN(n929) );
  NAND2_X4 U811 ( .A1(n2012), .A2(n2021), .ZN(n930) );
  XNOR2_X2 U812 ( .A(n585), .B(n936), .ZN(product[10]) );
  AOI21_X4 U813 ( .B1(n936), .B2(n932), .A(n933), .ZN(n931) );
  NAND2_X4 U816 ( .A1(n932), .A2(n935), .ZN(n585) );
  NOR2_X4 U818 ( .A1(n2022), .A2(n2029), .ZN(n934) );
  NAND2_X4 U819 ( .A1(n2022), .A2(n2029), .ZN(n935) );
  XNOR2_X2 U820 ( .A(n586), .B(n942), .ZN(product[9]) );
  AOI21_X4 U822 ( .B1(n942), .B2(n938), .A(n939), .ZN(n937) );
  NAND2_X4 U825 ( .A1(n938), .A2(n941), .ZN(n586) );
  NOR2_X4 U827 ( .A1(n2030), .A2(n2037), .ZN(n940) );
  NAND2_X4 U828 ( .A1(n2030), .A2(n2037), .ZN(n941) );
  XOR2_X2 U829 ( .A(n949), .B(n587), .Z(product[8]) );
  OAI21_X4 U830 ( .B1(n943), .B2(n955), .A(n944), .ZN(n942) );
  NAND2_X4 U831 ( .A1(n945), .A2(n950), .ZN(n943) );
  AOI21_X4 U832 ( .B1(n945), .B2(n951), .A(n946), .ZN(n944) );
  NAND2_X4 U835 ( .A1(n945), .A2(n948), .ZN(n587) );
  NOR2_X4 U837 ( .A1(n2038), .A2(n2043), .ZN(n947) );
  NAND2_X4 U838 ( .A1(n2038), .A2(n2043), .ZN(n948) );
  XNOR2_X2 U839 ( .A(n954), .B(n588), .ZN(product[7]) );
  AOI21_X4 U840 ( .B1(n954), .B2(n950), .A(n951), .ZN(n949) );
  NAND2_X4 U843 ( .A1(n950), .A2(n953), .ZN(n588) );
  NOR2_X4 U845 ( .A1(n2044), .A2(n2049), .ZN(n952) );
  NAND2_X4 U846 ( .A1(n2044), .A2(n2049), .ZN(n953) );
  XNOR2_X2 U847 ( .A(n589), .B(n960), .ZN(product[6]) );
  AOI21_X4 U849 ( .B1(n956), .B2(n960), .A(n957), .ZN(n955) );
  NAND2_X4 U852 ( .A1(n956), .A2(n959), .ZN(n589) );
  NOR2_X4 U854 ( .A1(n2050), .A2(n2053), .ZN(n958) );
  NAND2_X4 U855 ( .A1(n2050), .A2(n2053), .ZN(n959) );
  XOR2_X2 U856 ( .A(n590), .B(n963), .Z(product[5]) );
  OAI21_X4 U857 ( .B1(n961), .B2(n963), .A(n962), .ZN(n960) );
  NAND2_X4 U858 ( .A1(n1036), .A2(n962), .ZN(n590) );
  NOR2_X4 U860 ( .A1(n2054), .A2(n2057), .ZN(n961) );
  NAND2_X4 U861 ( .A1(n2054), .A2(n2057), .ZN(n962) );
  XNOR2_X2 U862 ( .A(n591), .B(n968), .ZN(product[4]) );
  AOI21_X4 U863 ( .B1(n964), .B2(n968), .A(n965), .ZN(n963) );
  NAND2_X4 U866 ( .A1(n964), .A2(n967), .ZN(n591) );
  NOR2_X4 U868 ( .A1(n2058), .A2(n2059), .ZN(n966) );
  NAND2_X4 U869 ( .A1(n2058), .A2(n2059), .ZN(n967) );
  XOR2_X2 U870 ( .A(n592), .B(n971), .Z(product[3]) );
  OAI21_X4 U871 ( .B1(n969), .B2(n971), .A(n970), .ZN(n968) );
  NAND2_X4 U872 ( .A1(n1038), .A2(n970), .ZN(n592) );
  NOR2_X4 U874 ( .A1(n2060), .A2(n2075), .ZN(n969) );
  NAND2_X4 U875 ( .A1(n2060), .A2(n2075), .ZN(n970) );
  XNOR2_X2 U876 ( .A(n593), .B(n976), .ZN(product[2]) );
  AOI21_X4 U877 ( .B1(n972), .B2(n976), .A(n973), .ZN(n971) );
  NAND2_X4 U880 ( .A1(n972), .A2(n975), .ZN(n593) );
  NOR2_X4 U882 ( .A1(n2603), .A2(n2635), .ZN(n974) );
  NAND2_X4 U883 ( .A1(n2603), .A2(n2635), .ZN(n975) );
  NAND2_X4 U886 ( .A1(n1040), .A2(n978), .ZN(n594) );
  NOR2_X4 U888 ( .A1(n2636), .A2(n2076), .ZN(n977) );
  NAND2_X4 U889 ( .A1(n2636), .A2(n2076), .ZN(n978) );
  FA_X1 U890 ( .A(n2095), .B(n1045), .CI(n1048), .CO(n1042), .S(n1043) );
  FA_X1 U892 ( .A(n1052), .B(n2128), .CI(n1049), .CO(n1046), .S(n1047) );
  FA_X1 U893 ( .A(n2078), .B(n1054), .CI(n2096), .CO(n1048), .S(n1049) );
  FA_X1 U894 ( .A(n1053), .B(n1060), .CI(n1058), .CO(n1050), .S(n1051) );
  FA_X1 U895 ( .A(n2129), .B(n1055), .CI(n2097), .CO(n1052), .S(n1053) );
  FA_X1 U897 ( .A(n1064), .B(n1061), .CI(n1059), .CO(n1056), .S(n1057) );
  FA_X1 U898 ( .A(n2162), .B(n2098), .CI(n1066), .CO(n1058), .S(n1059) );
  FA_X1 U899 ( .A(n2079), .B(n1068), .CI(n2130), .CO(n1060), .S(n1061) );
  FA_X1 U900 ( .A(n1072), .B(n1067), .CI(n1065), .CO(n1062), .S(n1063) );
  FA_X1 U901 ( .A(n1076), .B(n2099), .CI(n1074), .CO(n1064), .S(n1065) );
  FA_X1 U902 ( .A(n2163), .B(n1069), .CI(n2131), .CO(n1066), .S(n1067) );
  FA_X1 U904 ( .A(n1080), .B(n1082), .CI(n1073), .CO(n1070), .S(n1071) );
  FA_X1 U905 ( .A(n1077), .B(n1084), .CI(n1075), .CO(n1072), .S(n1073) );
  FA_X1 U906 ( .A(n2132), .B(n2100), .CI(n2196), .CO(n1074), .S(n1075) );
  FA_X1 U907 ( .A(n2080), .B(n1086), .CI(n2164), .CO(n1076), .S(n1077) );
  FA_X1 U908 ( .A(n1090), .B(n1083), .CI(n1081), .CO(n1078), .S(n1079) );
  FA_X1 U909 ( .A(n1085), .B(n1094), .CI(n1092), .CO(n1080), .S(n1081) );
  FA_X1 U910 ( .A(n2101), .B(n2133), .CI(n1096), .CO(n1082), .S(n1083) );
  FA_X1 U911 ( .A(n2197), .B(n1087), .CI(n2165), .CO(n1084), .S(n1085) );
  FA_X1 U913 ( .A(n1100), .B(n1093), .CI(n1091), .CO(n1088), .S(n1089) );
  FA_X1 U914 ( .A(n1095), .B(n1097), .CI(n1102), .CO(n1090), .S(n1091) );
  FA_X1 U915 ( .A(n1106), .B(n2230), .CI(n1104), .CO(n1092), .S(n1093) );
  FA_X1 U916 ( .A(n2102), .B(n2134), .CI(n2198), .CO(n1094), .S(n1095) );
  FA_X1 U917 ( .A(n2081), .B(n1108), .CI(n2166), .CO(n1096), .S(n1097) );
  FA_X1 U918 ( .A(n1112), .B(n1103), .CI(n1101), .CO(n1098), .S(n1099) );
  FA_X1 U919 ( .A(n1116), .B(n1105), .CI(n1114), .CO(n1100), .S(n1101) );
  FA_X1 U920 ( .A(n1118), .B(n1120), .CI(n1107), .CO(n1102), .S(n1103) );
  FA_X1 U921 ( .A(n2135), .B(n2103), .CI(n2167), .CO(n1104), .S(n1105) );
  FA_X1 U922 ( .A(n2231), .B(n1109), .CI(n2199), .CO(n1106), .S(n1107) );
  FA_X1 U924 ( .A(n1124), .B(n1115), .CI(n1113), .CO(n1110), .S(n1111) );
  FA_X1 U925 ( .A(n1117), .B(n1128), .CI(n1126), .CO(n1112), .S(n1113) );
  FA_X1 U926 ( .A(n1121), .B(n1130), .CI(n1119), .CO(n1114), .S(n1115) );
  FA_X1 U927 ( .A(n2264), .B(n2136), .CI(n1132), .CO(n1116), .S(n1117) );
  FA_X1 U928 ( .A(n2104), .B(n2168), .CI(n2232), .CO(n1118), .S(n1119) );
  FA_X1 U929 ( .A(n2082), .B(n1134), .CI(n2200), .CO(n1120), .S(n1121) );
  FA_X1 U930 ( .A(n1138), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U931 ( .A(n1129), .B(n1142), .CI(n1140), .CO(n1124), .S(n1125) );
  FA_X1 U932 ( .A(n1133), .B(n1144), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U933 ( .A(n1148), .B(n2137), .CI(n1146), .CO(n1128), .S(n1129) );
  FA_X1 U934 ( .A(n2105), .B(n2201), .CI(n2169), .CO(n1130), .S(n1131) );
  FA_X1 U935 ( .A(n2265), .B(n1135), .CI(n2233), .CO(n1132), .S(n1133) );
  FA_X1 U937 ( .A(n1152), .B(n1141), .CI(n1139), .CO(n1136), .S(n1137) );
  FA_X1 U938 ( .A(n1143), .B(n1156), .CI(n1154), .CO(n1138), .S(n1139) );
  FA_X1 U939 ( .A(n1145), .B(n1147), .CI(n1158), .CO(n1140), .S(n1141) );
  FA_X1 U940 ( .A(n1160), .B(n1162), .CI(n1149), .CO(n1142), .S(n1143) );
  FA_X1 U941 ( .A(n2266), .B(n2106), .CI(n2298), .CO(n1144), .S(n1145) );
  FA_X1 U942 ( .A(n2138), .B(n2170), .CI(n2234), .CO(n1146), .S(n1147) );
  FA_X1 U943 ( .A(n2083), .B(n1164), .CI(n2202), .CO(n1148), .S(n1149) );
  FA_X1 U944 ( .A(n1168), .B(n1155), .CI(n1153), .CO(n1150), .S(n1151) );
  FA_X1 U945 ( .A(n1157), .B(n1172), .CI(n1170), .CO(n1152), .S(n1153) );
  FA_X1 U946 ( .A(n1174), .B(n1161), .CI(n1159), .CO(n1154), .S(n1155) );
  FA_X1 U947 ( .A(n1176), .B(n1178), .CI(n1163), .CO(n1156), .S(n1157) );
  FA_X1 U948 ( .A(n2171), .B(n2203), .CI(n1180), .CO(n1158), .S(n1159) );
  FA_X1 U949 ( .A(n2107), .B(n2235), .CI(n2139), .CO(n1160), .S(n1161) );
  FA_X1 U950 ( .A(n2299), .B(n1165), .CI(n2267), .CO(n1162), .S(n1163) );
  FA_X1 U952 ( .A(n1184), .B(n1171), .CI(n1169), .CO(n1166), .S(n1167) );
  FA_X1 U953 ( .A(n1173), .B(n1188), .CI(n1186), .CO(n1168), .S(n1169) );
  FA_X1 U954 ( .A(n1190), .B(n1179), .CI(n1175), .CO(n1170), .S(n1171) );
  FA_X1 U955 ( .A(n1181), .B(n1192), .CI(n1177), .CO(n1172), .S(n1173) );
  FA_X1 U956 ( .A(n1196), .B(n2332), .CI(n1194), .CO(n1174), .S(n1175) );
  FA_X1 U957 ( .A(n2268), .B(n2140), .CI(n2300), .CO(n1176), .S(n1177) );
  FA_X1 U958 ( .A(n2108), .B(n2204), .CI(n2172), .CO(n1178), .S(n1179) );
  FA_X1 U959 ( .A(n2084), .B(n1198), .CI(n2236), .CO(n1180), .S(n1181) );
  FA_X1 U960 ( .A(n1202), .B(n1187), .CI(n1185), .CO(n1182), .S(n1183) );
  FA_X1 U961 ( .A(n1189), .B(n1206), .CI(n1204), .CO(n1184), .S(n1185) );
  FA_X1 U962 ( .A(n1208), .B(n1210), .CI(n1191), .CO(n1186), .S(n1187) );
  FA_X1 U963 ( .A(n1193), .B(n1197), .CI(n1195), .CO(n1188), .S(n1189) );
  FA_X1 U964 ( .A(n1214), .B(n1216), .CI(n1212), .CO(n1190), .S(n1191) );
  FA_X1 U965 ( .A(n2141), .B(n2205), .CI(n2173), .CO(n1192), .S(n1193) );
  FA_X1 U966 ( .A(n2109), .B(n2269), .CI(n2237), .CO(n1194), .S(n1195) );
  FA_X1 U967 ( .A(n2333), .B(n1199), .CI(n2301), .CO(n1196), .S(n1197) );
  FA_X1 U969 ( .A(n1220), .B(n1205), .CI(n1203), .CO(n1200), .S(n1201) );
  FA_X1 U970 ( .A(n1207), .B(n1224), .CI(n1222), .CO(n1202), .S(n1203) );
  FA_X1 U971 ( .A(n1211), .B(n1226), .CI(n1209), .CO(n1204), .S(n1205) );
  FA_X1 U972 ( .A(n1215), .B(n1213), .CI(n1228), .CO(n1206), .S(n1207) );
  FA_X1 U973 ( .A(n1230), .B(n1232), .CI(n1217), .CO(n1208), .S(n1209) );
  FA_X1 U974 ( .A(n2366), .B(n2334), .CI(n1234), .CO(n1210), .S(n1211) );
  FA_X1 U975 ( .A(n2302), .B(n2174), .CI(n2270), .CO(n1212), .S(n1213) );
  FA_X1 U976 ( .A(n2142), .B(n2206), .CI(n2110), .CO(n1214), .S(n1215) );
  FA_X1 U977 ( .A(n2085), .B(n1236), .CI(n2238), .CO(n1216), .S(n1217) );
  FA_X1 U978 ( .A(n1240), .B(n1223), .CI(n1221), .CO(n1218), .S(n1219) );
  FA_X1 U979 ( .A(n1225), .B(n1244), .CI(n1242), .CO(n1220), .S(n1221) );
  FA_X1 U980 ( .A(n1246), .B(n1229), .CI(n1227), .CO(n1222), .S(n1223) );
  FA_X1 U981 ( .A(n1233), .B(n1231), .CI(n1248), .CO(n1224), .S(n1225) );
  FA_X1 U982 ( .A(n1250), .B(n1252), .CI(n1235), .CO(n1226), .S(n1227) );
  FA_X1 U983 ( .A(n1256), .B(n2239), .CI(n1254), .CO(n1228), .S(n1229) );
  FA_X1 U984 ( .A(n2175), .B(n2271), .CI(n2207), .CO(n1230), .S(n1231) );
  FA_X1 U985 ( .A(n2111), .B(n2303), .CI(n2143), .CO(n1232), .S(n1233) );
  FA_X1 U986 ( .A(n2367), .B(n1237), .CI(n2335), .CO(n1234), .S(n1235) );
  FA_X1 U988 ( .A(n1260), .B(n1243), .CI(n1241), .CO(n1238), .S(n1239) );
  FA_X1 U989 ( .A(n1245), .B(n1264), .CI(n1262), .CO(n1240), .S(n1241) );
  FA_X1 U990 ( .A(n1249), .B(n1266), .CI(n1247), .CO(n1242), .S(n1243) );
  FA_X1 U991 ( .A(n1270), .B(n1251), .CI(n1268), .CO(n1244), .S(n1245) );
  FA_X1 U992 ( .A(n1253), .B(n1257), .CI(n1255), .CO(n1246), .S(n1247) );
  FA_X1 U993 ( .A(n1272), .B(n1276), .CI(n1274), .CO(n1248), .S(n1249) );
  FA_X1 U994 ( .A(n2336), .B(n2368), .CI(n2400), .CO(n1250), .S(n1251) );
  FA_X1 U995 ( .A(n2304), .B(n2144), .CI(n2208), .CO(n1252), .S(n1253) );
  FA_X1 U996 ( .A(n2112), .B(n2240), .CI(n2176), .CO(n1254), .S(n1255) );
  FA_X1 U997 ( .A(n2086), .B(n1278), .CI(n2272), .CO(n1256), .S(n1257) );
  FA_X1 U998 ( .A(n1282), .B(n1263), .CI(n1261), .CO(n1258), .S(n1259) );
  FA_X1 U999 ( .A(n1265), .B(n1286), .CI(n1284), .CO(n1260), .S(n1261) );
  FA_X1 U1000 ( .A(n1269), .B(n1288), .CI(n1267), .CO(n1262), .S(n1263) );
  FA_X1 U1001 ( .A(n1271), .B(n1292), .CI(n1290), .CO(n1264), .S(n1265) );
  FA_X1 U1002 ( .A(n1273), .B(n1277), .CI(n1275), .CO(n1266), .S(n1267) );
  FA_X1 U1003 ( .A(n1294), .B(n1298), .CI(n1296), .CO(n1268), .S(n1269) );
  FA_X1 U1004 ( .A(n2273), .B(n2305), .CI(n1300), .CO(n1270), .S(n1271) );
  FA_X1 U1005 ( .A(n2177), .B(n2241), .CI(n2209), .CO(n1272), .S(n1273) );
  FA_X1 U1006 ( .A(n2113), .B(n2337), .CI(n2145), .CO(n1274), .S(n1275) );
  FA_X1 U1007 ( .A(n2401), .B(n1279), .CI(n2369), .CO(n1276), .S(n1277) );
  FA_X1 U1011 ( .A(n1310), .B(n1291), .CI(n1289), .CO(n1284), .S(n1285) );
  FA_X1 U1012 ( .A(n1312), .B(n1314), .CI(n1293), .CO(n1286), .S(n1287) );
  FA_X1 U1013 ( .A(n1299), .B(n1295), .CI(n1297), .CO(n1288), .S(n1289) );
  FA_X1 U1014 ( .A(n1316), .B(n1318), .CI(n1301), .CO(n1290), .S(n1291) );
  FA_X1 U1015 ( .A(n1322), .B(n2434), .CI(n1320), .CO(n1292), .S(n1293) );
  FA_X1 U1016 ( .A(n2210), .B(n2402), .CI(n2370), .CO(n1294), .S(n1295) );
  FA_X1 U1017 ( .A(n2178), .B(n2306), .CI(n2338), .CO(n1296), .S(n1297) );
  FA_X1 U1018 ( .A(n2114), .B(n2242), .CI(n2146), .CO(n1298), .S(n1299) );
  FA_X1 U1019 ( .A(n2087), .B(n1324), .CI(n2274), .CO(n1300), .S(n1301) );
  FA_X1 U1020 ( .A(n1328), .B(n1307), .CI(n1305), .CO(n1302), .S(n1303) );
  FA_X1 U1021 ( .A(n1309), .B(n1332), .CI(n1330), .CO(n1304), .S(n1305) );
  FA_X1 U1022 ( .A(n1334), .B(n1313), .CI(n1311), .CO(n1306), .S(n1307) );
  FA_X1 U1023 ( .A(n1315), .B(n1338), .CI(n1336), .CO(n1308), .S(n1309) );
  FA_X1 U1024 ( .A(n1321), .B(n1319), .CI(n1340), .CO(n1310), .S(n1311) );
  FA_X1 U1025 ( .A(n1323), .B(n1342), .CI(n1317), .CO(n1312), .S(n1313) );
  FA_X1 U1026 ( .A(n1346), .B(n1348), .CI(n1344), .CO(n1314), .S(n1315) );
  FA_X1 U1027 ( .A(n2243), .B(n2307), .CI(n2275), .CO(n1316), .S(n1317) );
  FA_X1 U1028 ( .A(n2339), .B(n2179), .CI(n2211), .CO(n1318), .S(n1319) );
  FA_X1 U1029 ( .A(n2115), .B(n2371), .CI(n2147), .CO(n1320), .S(n1321) );
  FA_X1 U1030 ( .A(n2435), .B(n1325), .CI(n2403), .CO(n1322), .S(n1323) );
  FA_X1 U1032 ( .A(n1352), .B(n1331), .CI(n1329), .CO(n1326), .S(n1327) );
  FA_X1 U1033 ( .A(n1333), .B(n1356), .CI(n1354), .CO(n1328), .S(n1329) );
  FA_X1 U1034 ( .A(n1358), .B(n1337), .CI(n1335), .CO(n1330), .S(n1331) );
  FA_X1 U1035 ( .A(n1360), .B(n1341), .CI(n1339), .CO(n1332), .S(n1333) );
  FA_X1 U1036 ( .A(n1364), .B(n1347), .CI(n1362), .CO(n1334), .S(n1335) );
  FA_X1 U1037 ( .A(n1343), .B(n1349), .CI(n1345), .CO(n1336), .S(n1337) );
  FA_X1 U1038 ( .A(n1366), .B(n1370), .CI(n1368), .CO(n1338), .S(n1339) );
  FA_X1 U1039 ( .A(n2468), .B(n2436), .CI(n1372), .CO(n1340), .S(n1341) );
  FA_X1 U1040 ( .A(n2212), .B(n2404), .CI(n2372), .CO(n1342), .S(n1343) );
  FA_X1 U1041 ( .A(n2116), .B(n2340), .CI(n2244), .CO(n1344), .S(n1345) );
  FA_X1 U1042 ( .A(n2148), .B(n2276), .CI(n2180), .CO(n1346), .S(n1347) );
  FA_X1 U1043 ( .A(n2088), .B(n1374), .CI(n2308), .CO(n1348), .S(n1349) );
  FA_X1 U1044 ( .A(n1378), .B(n1355), .CI(n1353), .CO(n1350), .S(n1351) );
  FA_X1 U1045 ( .A(n1357), .B(n1382), .CI(n1380), .CO(n1352), .S(n1353) );
  FA_X1 U1046 ( .A(n1384), .B(n1361), .CI(n1359), .CO(n1354), .S(n1355) );
  FA_X1 U1047 ( .A(n1386), .B(n1365), .CI(n1363), .CO(n1356), .S(n1357) );
  FA_X1 U1048 ( .A(n1390), .B(n1369), .CI(n1388), .CO(n1358), .S(n1359) );
  FA_X1 U1049 ( .A(n1367), .B(n1373), .CI(n1371), .CO(n1360), .S(n1361) );
  FA_X1 U1050 ( .A(n1394), .B(n1396), .CI(n1392), .CO(n1362), .S(n1363) );
  FA_X1 U1051 ( .A(n1400), .B(n2341), .CI(n1398), .CO(n1364), .S(n1365) );
  FA_X1 U1052 ( .A(n2245), .B(n2373), .CI(n2309), .CO(n1366), .S(n1367) );
  FA_X1 U1053 ( .A(n2181), .B(n2405), .CI(n2213), .CO(n1368), .S(n1369) );
  FA_X1 U1054 ( .A(n2117), .B(n2437), .CI(n2149), .CO(n1370), .S(n1371) );
  FA_X1 U1055 ( .A(n2469), .B(n1375), .CI(n2277), .CO(n1372), .S(n1373) );
  FA_X1 U1058 ( .A(n1383), .B(n1408), .CI(n1406), .CO(n1378), .S(n1379) );
  FA_X1 U1059 ( .A(n1410), .B(n1387), .CI(n1385), .CO(n1380), .S(n1381) );
  FA_X1 U1060 ( .A(n1389), .B(n1391), .CI(n1412), .CO(n1382), .S(n1383) );
  FA_X1 U1061 ( .A(n1416), .B(n1418), .CI(n1414), .CO(n1384), .S(n1385) );
  FA_X1 U1062 ( .A(n1399), .B(n1397), .CI(n1393), .CO(n1386), .S(n1387) );
  FA_X1 U1063 ( .A(n1401), .B(n1422), .CI(n1395), .CO(n1388), .S(n1389) );
  FA_X1 U1064 ( .A(n1420), .B(n1426), .CI(n1424), .CO(n1390), .S(n1391) );
  FA_X1 U1065 ( .A(n2438), .B(n2470), .CI(n2502), .CO(n1392), .S(n1393) );
  FA_X1 U1066 ( .A(n2374), .B(n2246), .CI(n2406), .CO(n1394), .S(n1395) );
  FA_X1 U1067 ( .A(n2214), .B(n2310), .CI(n2118), .CO(n1396), .S(n1397) );
  FA_X1 U1068 ( .A(n2150), .B(n2182), .CI(n2278), .CO(n1398), .S(n1399) );
  FA_X1 U1069 ( .A(n2089), .B(n1428), .CI(n2342), .CO(n1400), .S(n1401) );
  FA_X1 U1071 ( .A(n1409), .B(n1436), .CI(n1434), .CO(n1404), .S(n1405) );
  FA_X1 U1072 ( .A(n1438), .B(n1413), .CI(n1411), .CO(n1406), .S(n1407) );
  FA_X1 U1073 ( .A(n1415), .B(n1417), .CI(n1440), .CO(n1408), .S(n1409) );
  FA_X1 U1074 ( .A(n1419), .B(n1444), .CI(n1442), .CO(n1410), .S(n1411) );
  FA_X1 U1075 ( .A(n1425), .B(n1423), .CI(n1446), .CO(n1412), .S(n1413) );
  FA_X1 U1076 ( .A(n1427), .B(n1452), .CI(n1421), .CO(n1414), .S(n1415) );
  FA_X1 U1077 ( .A(n1448), .B(n1454), .CI(n1450), .CO(n1416), .S(n1417) );
  FA_X1 U1078 ( .A(n2247), .B(n2311), .CI(n1456), .CO(n1418), .S(n1419) );
  FA_X1 U1079 ( .A(n2183), .B(n2343), .CI(n2215), .CO(n1420), .S(n1421) );
  FA_X1 U1081 ( .A(n2439), .B(n2279), .CI(n2119), .CO(n1424), .S(n1425) );
  FA_X1 U1082 ( .A(n2503), .B(n1429), .CI(n2471), .CO(n1426), .S(n1427) );
  FA_X1 U1084 ( .A(n1460), .B(n1435), .CI(n1433), .CO(n1430), .S(n1431) );
  FA_X1 U1086 ( .A(n1466), .B(n1441), .CI(n1439), .CO(n1434), .S(n1435) );
  FA_X1 U1087 ( .A(n1443), .B(n1445), .CI(n1468), .CO(n1436), .S(n1437) );
  FA_X1 U1088 ( .A(n1472), .B(n1447), .CI(n1470), .CO(n1438), .S(n1439) );
  FA_X1 U1089 ( .A(n1453), .B(n1455), .CI(n1474), .CO(n1440), .S(n1441) );
  FA_X1 U1090 ( .A(n1449), .B(n1457), .CI(n1451), .CO(n1442), .S(n1443) );
  FA_X1 U1091 ( .A(n1482), .B(n1478), .CI(n1480), .CO(n1444), .S(n1445) );
  FA_X1 U1092 ( .A(n2536), .B(n1484), .CI(n1476), .CO(n1446), .S(n1447) );
  FA_X1 U1093 ( .A(n2504), .B(n2472), .CI(n2280), .CO(n1448), .S(n1449) );
  FA_X1 U1094 ( .A(n2408), .B(n2248), .CI(n2440), .CO(n1450), .S(n1451) );
  FA_X1 U1095 ( .A(n2152), .B(n2376), .CI(n2216), .CO(n1452), .S(n1453) );
  FA_X1 U1096 ( .A(n2120), .B(n2312), .CI(n2184), .CO(n1454), .S(n1455) );
  FA_X1 U1097 ( .A(n2090), .B(n1486), .CI(n2344), .CO(n1456), .S(n1457) );
  FA_X1 U1098 ( .A(n1490), .B(n1463), .CI(n1461), .CO(n1458), .S(n1459) );
  FA_X1 U1100 ( .A(n1496), .B(n1469), .CI(n1467), .CO(n1462), .S(n1463) );
  FA_X1 U1101 ( .A(n1471), .B(n1473), .CI(n1498), .CO(n1464), .S(n1465) );
  FA_X1 U1102 ( .A(n1475), .B(n1502), .CI(n1500), .CO(n1466), .S(n1467) );
  FA_X1 U1103 ( .A(n1506), .B(n1481), .CI(n1504), .CO(n1468), .S(n1469) );
  FA_X1 U1104 ( .A(n1483), .B(n1477), .CI(n1479), .CO(n1470), .S(n1471) );
  FA_X1 U1105 ( .A(n1514), .B(n1512), .CI(n1485), .CO(n1472), .S(n1473) );
  FA_X1 U1106 ( .A(n1508), .B(n1516), .CI(n1510), .CO(n1474), .S(n1475) );
  FA_X1 U1107 ( .A(n2249), .B(n2313), .CI(n2345), .CO(n1476), .S(n1477) );
  FA_X1 U1108 ( .A(n2185), .B(n2377), .CI(n2217), .CO(n1478), .S(n1479) );
  FA_X1 U1109 ( .A(n2153), .B(n2441), .CI(n2409), .CO(n1480), .S(n1481) );
  FA_X1 U1110 ( .A(n2473), .B(n2281), .CI(n2121), .CO(n1482), .S(n1483) );
  FA_X1 U1111 ( .A(n2505), .B(n1487), .CI(n2537), .CO(n1484), .S(n1485) );
  FA_X1 U1115 ( .A(n1499), .B(n1526), .CI(n1497), .CO(n1492), .S(n1493) );
  FA_X1 U1116 ( .A(n1501), .B(n1503), .CI(n1528), .CO(n1494), .S(n1495) );
  FA_X1 U1117 ( .A(n1505), .B(n1532), .CI(n1530), .CO(n1496), .S(n1497) );
  FA_X1 U1118 ( .A(n1534), .B(n1536), .CI(n1507), .CO(n1498), .S(n1499) );
  FA_X1 U1119 ( .A(n1515), .B(n1513), .CI(n1511), .CO(n1500), .S(n1501) );
  FA_X1 U1120 ( .A(n1517), .B(n1540), .CI(n1509), .CO(n1502), .S(n1503) );
  FA_X1 U1121 ( .A(n1544), .B(n1538), .CI(n1542), .CO(n1504), .S(n1505) );
  FA_X1 U1122 ( .A(n2570), .B(n2474), .CI(n1546), .CO(n1506), .S(n1507) );
  FA_X1 U1123 ( .A(n2506), .B(n2538), .CI(n2442), .CO(n1508), .S(n1509) );
  FA_X1 U1124 ( .A(n2346), .B(n2250), .CI(n2282), .CO(n1510), .S(n1511) );
  FA_X1 U1125 ( .A(n2218), .B(n2410), .CI(n2186), .CO(n1512), .S(n1513) );
  FA_X1 U1126 ( .A(n2122), .B(n2314), .CI(n2154), .CO(n1514), .S(n1515) );
  FA_X1 U1127 ( .A(n2091), .B(n1548), .CI(n2378), .CO(n1516), .S(n1517) );
  FA_X1 U1130 ( .A(n1529), .B(n1558), .CI(n1527), .CO(n1522), .S(n1523) );
  FA_X1 U1131 ( .A(n1531), .B(n1533), .CI(n1560), .CO(n1524), .S(n1525) );
  FA_X1 U1132 ( .A(n1562), .B(n1537), .CI(n1535), .CO(n1526), .S(n1527) );
  FA_X1 U1133 ( .A(n1566), .B(n1568), .CI(n1564), .CO(n1528), .S(n1529) );
  FA_X1 U1134 ( .A(n1545), .B(n1543), .CI(n1541), .CO(n1530), .S(n1531) );
  FA_X1 U1135 ( .A(n1547), .B(n1572), .CI(n1539), .CO(n1532), .S(n1533) );
  FA_X1 U1136 ( .A(n1576), .B(n1570), .CI(n1574), .CO(n1534), .S(n1535) );
  FA_X1 U1137 ( .A(n2411), .B(n2379), .CI(n1578), .CO(n1536), .S(n1537) );
  FA_X1 U1138 ( .A(n2315), .B(n2347), .CI(n2443), .CO(n1538), .S(n1539) );
  FA_X1 U1139 ( .A(n2475), .B(n2251), .CI(n2283), .CO(n1540), .S(n1541) );
  FA_X1 U1140 ( .A(n2187), .B(n2507), .CI(n2219), .CO(n1542), .S(n1543) );
  FA_X1 U1142 ( .A(n1580), .B(n2092), .CI(n2571), .CO(n1546), .S(n1547) );
  FA_X1 U1145 ( .A(n1557), .B(n1559), .CI(n1585), .CO(n1552), .S(n1553) );
  FA_X1 U1146 ( .A(n1561), .B(n1589), .CI(n1587), .CO(n1554), .S(n1555) );
  FA_X1 U1147 ( .A(n1591), .B(n1565), .CI(n1563), .CO(n1556), .S(n1557) );
  FA_X1 U1148 ( .A(n1593), .B(n1569), .CI(n1567), .CO(n1558), .S(n1559) );
  FA_X1 U1149 ( .A(n1597), .B(n1575), .CI(n1595), .CO(n1560), .S(n1561) );
  FA_X1 U1151 ( .A(n1599), .B(n1605), .CI(n1579), .CO(n1564), .S(n1565) );
  FA_X1 U1152 ( .A(n1607), .B(n1601), .CI(n1603), .CO(n1566), .S(n1567) );
  FA_X1 U1153 ( .A(n2604), .B(n2508), .CI(n1609), .CO(n1568), .S(n1569) );
  FA_X1 U1154 ( .A(n2476), .B(n2540), .CI(n2572), .CO(n1570), .S(n1571) );
  FA_X1 U1155 ( .A(n2284), .B(n2380), .CI(n2316), .CO(n1572), .S(n1573) );
  FA_X1 U1156 ( .A(n2252), .B(n2444), .CI(n2220), .CO(n1574), .S(n1575) );
  FA_X1 U1158 ( .A(n2412), .B(n1580), .CI(n2156), .CO(n1578), .S(n1579) );
  FA_X1 U1160 ( .A(n1613), .B(n1586), .CI(n1584), .CO(n1581), .S(n1582) );
  FA_X1 U1161 ( .A(n1588), .B(n1590), .CI(n1615), .CO(n1583), .S(n1584) );
  FA_X1 U1162 ( .A(n1619), .B(n1592), .CI(n1617), .CO(n1585), .S(n1586) );
  FA_X1 U1163 ( .A(n1621), .B(n1596), .CI(n1594), .CO(n1587), .S(n1588) );
  FA_X1 U1164 ( .A(n1623), .B(n1625), .CI(n1598), .CO(n1589), .S(n1590) );
  FA_X1 U1165 ( .A(n1600), .B(n1606), .CI(n1627), .CO(n1591), .S(n1592) );
  FA_X1 U1166 ( .A(n1608), .B(n1602), .CI(n1604), .CO(n1593), .S(n1594) );
  FA_X1 U1167 ( .A(n1633), .B(n1629), .CI(n1610), .CO(n1595), .S(n1596) );
  FA_X1 U1168 ( .A(n1637), .B(n1631), .CI(n1635), .CO(n1597), .S(n1598) );
  FA_X1 U1169 ( .A(n2445), .B(n2413), .CI(n1639), .CO(n1599), .S(n1600) );
  FA_X1 U1170 ( .A(n2349), .B(n2477), .CI(n2317), .CO(n1601), .S(n1602) );
  FA_X1 U1171 ( .A(n2253), .B(n2509), .CI(n2285), .CO(n1603), .S(n1604) );
  FA_X1 U1172 ( .A(n2541), .B(n2381), .CI(n2221), .CO(n1605), .S(n1606) );
  FA_X1 U1173 ( .A(n2125), .B(n2573), .CI(n2189), .CO(n1607), .S(n1608) );
  FA_X1 U1174 ( .A(n2157), .B(n2093), .CI(n2605), .CO(n1609), .S(n1610) );
  FA_X1 U1175 ( .A(n1643), .B(n1616), .CI(n1614), .CO(n1611), .S(n1612) );
  FA_X1 U1176 ( .A(n1618), .B(n1620), .CI(n1645), .CO(n1613), .S(n1614) );
  FA_X1 U1177 ( .A(n1649), .B(n1622), .CI(n1647), .CO(n1615), .S(n1616) );
  FA_X1 U1178 ( .A(n1651), .B(n1626), .CI(n1624), .CO(n1617), .S(n1618) );
  FA_X1 U1179 ( .A(n1628), .B(n1655), .CI(n1653), .CO(n1619), .S(n1620) );
  FA_X1 U1180 ( .A(n1632), .B(n1634), .CI(n1657), .CO(n1621), .S(n1622) );
  FA_X1 U1181 ( .A(n1638), .B(n1630), .CI(n1636), .CO(n1623), .S(n1624) );
  FA_X1 U1182 ( .A(n1663), .B(n1659), .CI(n1661), .CO(n1625), .S(n1626) );
  FA_X1 U1183 ( .A(n1667), .B(n1640), .CI(n1665), .CO(n1627), .S(n1628) );
  FA_X1 U1184 ( .A(n2414), .B(n2286), .CI(n2350), .CO(n1629), .S(n1630) );
  FA_X1 U1185 ( .A(n2190), .B(n2446), .CI(n2222), .CO(n1631), .S(n1632) );
  FA_X1 U1186 ( .A(n2158), .B(n2254), .CI(n2478), .CO(n1633), .S(n1634) );
  FA_X1 U1187 ( .A(n2542), .B(n2318), .CI(n2510), .CO(n1635), .S(n1636) );
  FA_X1 U1188 ( .A(n2606), .B(n2382), .CI(n2574), .CO(n1637), .S(n1638) );
  HA_X1 U1189 ( .A(n2126), .B(n2061), .CO(n1639), .S(n1640) );
  FA_X1 U1191 ( .A(n1648), .B(n1650), .CI(n1673), .CO(n1643), .S(n1644) );
  FA_X1 U1192 ( .A(n1677), .B(n1652), .CI(n1675), .CO(n1645), .S(n1646) );
  FA_X1 U1193 ( .A(n1656), .B(n1679), .CI(n1654), .CO(n1647), .S(n1648) );
  FA_X1 U1194 ( .A(n1681), .B(n1683), .CI(n1658), .CO(n1649), .S(n1650) );
  FA_X1 U1195 ( .A(n1664), .B(n1662), .CI(n1685), .CO(n1651), .S(n1652) );
  FA_X1 U1196 ( .A(n1668), .B(n1660), .CI(n1666), .CO(n1653), .S(n1654) );
  FA_X1 U1197 ( .A(n1691), .B(n1687), .CI(n1689), .CO(n1655), .S(n1656) );
  FA_X1 U1198 ( .A(n1695), .B(n2447), .CI(n1693), .CO(n1657), .S(n1658) );
  FA_X1 U1199 ( .A(n2383), .B(n2479), .CI(n2415), .CO(n1659), .S(n1660) );
  FA_X1 U1200 ( .A(n2319), .B(n2287), .CI(n2351), .CO(n1661), .S(n1662) );
  FA_X1 U1201 ( .A(n2223), .B(n2511), .CI(n2255), .CO(n1663), .S(n1664) );
  FA_X1 U1202 ( .A(n2191), .B(n2543), .CI(n2575), .CO(n1665), .S(n1666) );
  FA_X1 U1204 ( .A(n1699), .B(n1674), .CI(n1672), .CO(n1669), .S(n1670) );
  FA_X1 U1206 ( .A(n1705), .B(n1680), .CI(n1703), .CO(n1673), .S(n1674) );
  FA_X1 U1207 ( .A(n1684), .B(n1707), .CI(n1682), .CO(n1675), .S(n1676) );
  FA_X1 U1208 ( .A(n1686), .B(n1711), .CI(n1709), .CO(n1677), .S(n1678) );
  FA_X1 U1209 ( .A(n1690), .B(n1692), .CI(n1694), .CO(n1679), .S(n1680) );
  FA_X1 U1210 ( .A(n1713), .B(n1717), .CI(n1688), .CO(n1681), .S(n1682) );
  FA_X1 U1211 ( .A(n1721), .B(n1715), .CI(n1719), .CO(n1683), .S(n1684) );
  FA_X1 U1212 ( .A(n2480), .B(n2448), .CI(n1696), .CO(n1685), .S(n1686) );
  FA_X1 U1213 ( .A(n2512), .B(n2320), .CI(n2288), .CO(n1687), .S(n1688) );
  FA_X1 U1214 ( .A(n2256), .B(n2416), .CI(n2544), .CO(n1689), .S(n1690) );
  FA_X1 U1215 ( .A(n2224), .B(n2352), .CI(n2576), .CO(n1691), .S(n1692) );
  FA_X1 U1216 ( .A(n2608), .B(n2384), .CI(n2192), .CO(n1693), .S(n1694) );
  HA_X1 U1217 ( .A(n2160), .B(n2062), .CO(n1695), .S(n1696) );
  FA_X1 U1218 ( .A(n1725), .B(n1702), .CI(n1700), .CO(n1697), .S(n1698) );
  FA_X1 U1219 ( .A(n1704), .B(n1729), .CI(n1727), .CO(n1699), .S(n1700) );
  FA_X1 U1220 ( .A(n1731), .B(n1708), .CI(n1706), .CO(n1701), .S(n1702) );
  FA_X1 U1221 ( .A(n1733), .B(n1712), .CI(n1710), .CO(n1703), .S(n1704) );
  FA_X1 U1222 ( .A(n1737), .B(n1718), .CI(n1735), .CO(n1705), .S(n1706) );
  FA_X1 U1223 ( .A(n1722), .B(n1716), .CI(n1720), .CO(n1707), .S(n1708) );
  FA_X1 U1224 ( .A(n1741), .B(n1739), .CI(n1714), .CO(n1709), .S(n1710) );
  FA_X1 U1225 ( .A(n1745), .B(n1747), .CI(n1743), .CO(n1711), .S(n1712) );
  FA_X1 U1226 ( .A(n2385), .B(n2417), .CI(n2449), .CO(n1713), .S(n1714) );
  FA_X1 U1227 ( .A(n2321), .B(n2481), .CI(n2353), .CO(n1715), .S(n1716) );
  FA_X1 U1228 ( .A(n2257), .B(n2513), .CI(n2289), .CO(n1717), .S(n1718) );
  FA_X1 U1229 ( .A(n2225), .B(n2577), .CI(n2545), .CO(n1719), .S(n1720) );
  FA_X1 U1230 ( .A(n2193), .B(n2609), .CI(n2161), .CO(n1721), .S(n1722) );
  FA_X1 U1231 ( .A(n1751), .B(n1728), .CI(n1726), .CO(n1723), .S(n1724) );
  FA_X1 U1232 ( .A(n1730), .B(n1732), .CI(n1753), .CO(n1725), .S(n1726) );
  FA_X1 U1233 ( .A(n1734), .B(n1757), .CI(n1755), .CO(n1727), .S(n1728) );
  FA_X1 U1235 ( .A(n1744), .B(n1746), .CI(n1761), .CO(n1731), .S(n1732) );
  FA_X1 U1236 ( .A(n1740), .B(n1763), .CI(n1742), .CO(n1733), .S(n1734) );
  FA_X1 U1237 ( .A(n1767), .B(n1765), .CI(n1769), .CO(n1735), .S(n1736) );
  FA_X1 U1238 ( .A(n1748), .B(n2514), .CI(n1771), .CO(n1737), .S(n1738) );
  FA_X1 U1239 ( .A(n2450), .B(n2546), .CI(n2482), .CO(n1739), .S(n1740) );
  FA_X1 U1240 ( .A(n2578), .B(n2354), .CI(n2322), .CO(n1741), .S(n1742) );
  FA_X1 U1241 ( .A(n2258), .B(n2386), .CI(n2290), .CO(n1743), .S(n1744) );
  FA_X1 U1242 ( .A(n2226), .B(n2418), .CI(n2610), .CO(n1745), .S(n1746) );
  HA_X1 U1243 ( .A(n2194), .B(n2063), .CO(n1747), .S(n1748) );
  FA_X1 U1244 ( .A(n1775), .B(n1754), .CI(n1752), .CO(n1749), .S(n1750) );
  FA_X1 U1245 ( .A(n1779), .B(n1777), .CI(n1756), .CO(n1751), .S(n1752) );
  FA_X1 U1246 ( .A(n1758), .B(n1762), .CI(n1760), .CO(n1753), .S(n1754) );
  FA_X1 U1247 ( .A(n1783), .B(n1785), .CI(n1781), .CO(n1755), .S(n1756) );
  FA_X1 U1248 ( .A(n1770), .B(n1772), .CI(n1764), .CO(n1757), .S(n1758) );
  FA_X1 U1249 ( .A(n1766), .B(n1793), .CI(n1768), .CO(n1759), .S(n1760) );
  FA_X1 U1250 ( .A(n1787), .B(n1789), .CI(n1791), .CO(n1761), .S(n1762) );
  FA_X1 U1251 ( .A(n2451), .B(n2483), .CI(n1795), .CO(n1763), .S(n1764) );
  FA_X1 U1252 ( .A(n2387), .B(n2515), .CI(n2419), .CO(n1765), .S(n1766) );
  FA_X1 U1253 ( .A(n2323), .B(n2547), .CI(n2355), .CO(n1767), .S(n1768) );
  FA_X1 U1254 ( .A(n2259), .B(n2579), .CI(n2291), .CO(n1769), .S(n1770) );
  FA_X1 U1255 ( .A(n2227), .B(n2611), .CI(n2195), .CO(n1771), .S(n1772) );
  FA_X1 U1256 ( .A(n1799), .B(n1778), .CI(n1776), .CO(n1773), .S(n1774) );
  FA_X1 U1257 ( .A(n1780), .B(n1803), .CI(n1801), .CO(n1775), .S(n1776) );
  FA_X1 U1258 ( .A(n1784), .B(n1805), .CI(n1782), .CO(n1777), .S(n1778) );
  FA_X1 U1259 ( .A(n1807), .B(n1809), .CI(n1786), .CO(n1779), .S(n1780) );
  FA_X1 U1260 ( .A(n1794), .B(n1790), .CI(n1792), .CO(n1781), .S(n1782) );
  FA_X1 U1261 ( .A(n1811), .B(n1813), .CI(n1788), .CO(n1783), .S(n1784) );
  FA_X1 U1262 ( .A(n1817), .B(n1796), .CI(n1815), .CO(n1785), .S(n1786) );
  FA_X1 U1263 ( .A(n2356), .B(n2484), .CI(n2452), .CO(n1787), .S(n1788) );
  FA_X1 U1264 ( .A(n2292), .B(n2516), .CI(n2324), .CO(n1789), .S(n1790) );
  FA_X1 U1265 ( .A(n2580), .B(n2388), .CI(n2548), .CO(n1791), .S(n1792) );
  FA_X1 U1266 ( .A(n2612), .B(n2420), .CI(n2260), .CO(n1793), .S(n1794) );
  HA_X1 U1267 ( .A(n2228), .B(n2064), .CO(n1795), .S(n1796) );
  FA_X1 U1268 ( .A(n1821), .B(n1802), .CI(n1800), .CO(n1797), .S(n1798) );
  FA_X1 U1269 ( .A(n1804), .B(n1825), .CI(n1823), .CO(n1799), .S(n1800) );
  FA_X1 U1270 ( .A(n1808), .B(n1827), .CI(n1806), .CO(n1801), .S(n1802) );
  FA_X1 U1271 ( .A(n1829), .B(n1831), .CI(n1810), .CO(n1803), .S(n1804) );
  FA_X1 U1272 ( .A(n1818), .B(n1814), .CI(n1816), .CO(n1805), .S(n1806) );
  FA_X1 U1273 ( .A(n1833), .B(n1835), .CI(n1812), .CO(n1807), .S(n1808) );
  FA_X1 U1274 ( .A(n1839), .B(n2453), .CI(n1837), .CO(n1809), .S(n1810) );
  FA_X1 U1275 ( .A(n2389), .B(n2485), .CI(n2421), .CO(n1811), .S(n1812) );
  FA_X1 U1276 ( .A(n2357), .B(n2549), .CI(n2517), .CO(n1813), .S(n1814) );
  FA_X1 U1277 ( .A(n2293), .B(n2581), .CI(n2325), .CO(n1815), .S(n1816) );
  FA_X1 U1278 ( .A(n2261), .B(n2613), .CI(n2229), .CO(n1817), .S(n1818) );
  FA_X1 U1279 ( .A(n1843), .B(n1824), .CI(n1822), .CO(n1819), .S(n1820) );
  FA_X1 U1280 ( .A(n1845), .B(n1828), .CI(n1826), .CO(n1821), .S(n1822) );
  FA_X1 U1281 ( .A(n1830), .B(n1849), .CI(n1847), .CO(n1823), .S(n1824) );
  FA_X1 U1282 ( .A(n1851), .B(n1838), .CI(n1832), .CO(n1825), .S(n1826) );
  FA_X1 U1283 ( .A(n1834), .B(n1857), .CI(n1836), .CO(n1827), .S(n1828) );
  FA_X1 U1284 ( .A(n1853), .B(n1859), .CI(n1855), .CO(n1829), .S(n1830) );
  FA_X1 U1285 ( .A(n2486), .B(n2518), .CI(n1840), .CO(n1831), .S(n1832) );
  FA_X1 U1286 ( .A(n2358), .B(n2550), .CI(n2390), .CO(n1833), .S(n1834) );
  FA_X1 U1287 ( .A(n2326), .B(n2422), .CI(n2582), .CO(n1835), .S(n1836) );
  FA_X1 U1288 ( .A(n2614), .B(n2454), .CI(n2294), .CO(n1837), .S(n1838) );
  HA_X1 U1289 ( .A(n2262), .B(n2065), .CO(n1839), .S(n1840) );
  FA_X1 U1290 ( .A(n1863), .B(n1846), .CI(n1844), .CO(n1841), .S(n1842) );
  FA_X1 U1291 ( .A(n1848), .B(n1850), .CI(n1865), .CO(n1843), .S(n1844) );
  FA_X1 U1292 ( .A(n1852), .B(n1869), .CI(n1867), .CO(n1845), .S(n1846) );
  FA_X1 U1293 ( .A(n1860), .B(n1858), .CI(n1871), .CO(n1847), .S(n1848) );
  FA_X1 U1294 ( .A(n1854), .B(n1873), .CI(n1856), .CO(n1849), .S(n1850) );
  FA_X1 U1295 ( .A(n1877), .B(n1879), .CI(n1875), .CO(n1851), .S(n1852) );
  FA_X1 U1296 ( .A(n2455), .B(n2519), .CI(n2487), .CO(n1853), .S(n1854) );
  FA_X1 U1297 ( .A(n2391), .B(n2551), .CI(n2423), .CO(n1855), .S(n1856) );
  FA_X1 U1298 ( .A(n2327), .B(n2583), .CI(n2359), .CO(n1857), .S(n1858) );
  FA_X1 U1299 ( .A(n2295), .B(n2615), .CI(n2263), .CO(n1859), .S(n1860) );
  FA_X1 U1300 ( .A(n1883), .B(n1866), .CI(n1864), .CO(n1861), .S(n1862) );
  FA_X1 U1301 ( .A(n1868), .B(n1870), .CI(n1885), .CO(n1863), .S(n1864) );
  FA_X1 U1302 ( .A(n1872), .B(n1889), .CI(n1887), .CO(n1865), .S(n1866) );
  FA_X1 U1303 ( .A(n1878), .B(n1874), .CI(n1876), .CO(n1867), .S(n1868) );
  FA_X1 U1304 ( .A(n1893), .B(n1895), .CI(n1891), .CO(n1869), .S(n1870) );
  FA_X1 U1305 ( .A(n1880), .B(n2488), .CI(n1897), .CO(n1871), .S(n1872) );
  FA_X1 U1306 ( .A(n2360), .B(n2392), .CI(n2520), .CO(n1873), .S(n1874) );
  FA_X1 U1307 ( .A(n2328), .B(n2424), .CI(n2552), .CO(n1875), .S(n1876) );
  FA_X1 U1308 ( .A(n2616), .B(n2584), .CI(n2456), .CO(n1877), .S(n1878) );
  HA_X1 U1309 ( .A(n2296), .B(n2066), .CO(n1879), .S(n1880) );
  FA_X1 U1310 ( .A(n1901), .B(n1886), .CI(n1884), .CO(n1881), .S(n1882) );
  FA_X1 U1311 ( .A(n1888), .B(n1890), .CI(n1903), .CO(n1883), .S(n1884) );
  FA_X1 U1312 ( .A(n1907), .B(n1892), .CI(n1905), .CO(n1885), .S(n1886) );
  FA_X1 U1313 ( .A(n1898), .B(n1894), .CI(n1896), .CO(n1887), .S(n1888) );
  FA_X1 U1314 ( .A(n1909), .B(n1913), .CI(n1911), .CO(n1889), .S(n1890) );
  FA_X1 U1315 ( .A(n2489), .B(n2521), .CI(n1915), .CO(n1891), .S(n1892) );
  FA_X1 U1316 ( .A(n2425), .B(n2553), .CI(n2457), .CO(n1893), .S(n1894) );
  FA_X1 U1317 ( .A(n2361), .B(n2585), .CI(n2393), .CO(n1895), .S(n1896) );
  FA_X1 U1318 ( .A(n2329), .B(n2617), .CI(n2297), .CO(n1897), .S(n1898) );
  FA_X1 U1319 ( .A(n1919), .B(n1904), .CI(n1902), .CO(n1899), .S(n1900) );
  FA_X1 U1320 ( .A(n1906), .B(n1923), .CI(n1921), .CO(n1901), .S(n1902) );
  FA_X1 U1321 ( .A(n1925), .B(n1914), .CI(n1908), .CO(n1903), .S(n1904) );
  FA_X1 U1322 ( .A(n1910), .B(n1927), .CI(n1912), .CO(n1905), .S(n1906) );
  FA_X1 U1323 ( .A(n1931), .B(n1916), .CI(n1929), .CO(n1907), .S(n1908) );
  FA_X1 U1324 ( .A(n2554), .B(n2586), .CI(n2458), .CO(n1909), .S(n1910) );
  FA_X1 U1325 ( .A(n2618), .B(n2522), .CI(n2426), .CO(n1911), .S(n1912) );
  FA_X1 U1326 ( .A(n2362), .B(n2490), .CI(n2394), .CO(n1913), .S(n1914) );
  HA_X1 U1327 ( .A(n2330), .B(n2067), .CO(n1915), .S(n1916) );
  FA_X1 U1329 ( .A(n1924), .B(n1926), .CI(n1937), .CO(n1919), .S(n1920) );
  FA_X1 U1330 ( .A(n1941), .B(n1932), .CI(n1939), .CO(n1921), .S(n1922) );
  FA_X1 U1331 ( .A(n1928), .B(n1943), .CI(n1930), .CO(n1923), .S(n1924) );
  FA_X1 U1332 ( .A(n1947), .B(n2523), .CI(n1945), .CO(n1925), .S(n1926) );
  FA_X1 U1333 ( .A(n2491), .B(n2555), .CI(n2459), .CO(n1927), .S(n1928) );
  FA_X1 U1334 ( .A(n2395), .B(n2587), .CI(n2427), .CO(n1929), .S(n1930) );
  FA_X1 U1335 ( .A(n2363), .B(n2619), .CI(n2331), .CO(n1931), .S(n1932) );
  FA_X1 U1336 ( .A(n1938), .B(n1951), .CI(n1936), .CO(n1933), .S(n1934) );
  FA_X1 U1337 ( .A(n1953), .B(n1942), .CI(n1940), .CO(n1935), .S(n1936) );
  FA_X1 U1338 ( .A(n1946), .B(n1944), .CI(n1955), .CO(n1937), .S(n1938) );
  FA_X1 U1339 ( .A(n1957), .B(n1961), .CI(n1959), .CO(n1939), .S(n1940) );
  FA_X1 U1340 ( .A(n2556), .B(n2588), .CI(n1948), .CO(n1941), .S(n1942) );
  FA_X1 U1341 ( .A(n2428), .B(n2524), .CI(n2460), .CO(n1943), .S(n1944) );
  FA_X1 U1342 ( .A(n2396), .B(n2492), .CI(n2620), .CO(n1945), .S(n1946) );
  HA_X1 U1343 ( .A(n2364), .B(n2068), .CO(n1947), .S(n1948) );
  FA_X1 U1344 ( .A(n1965), .B(n1954), .CI(n1952), .CO(n1949), .S(n1950) );
  FA_X1 U1345 ( .A(n1967), .B(n1969), .CI(n1956), .CO(n1951), .S(n1952) );
  FA_X1 U1346 ( .A(n1960), .B(n1962), .CI(n1958), .CO(n1953), .S(n1954) );
  FA_X1 U1347 ( .A(n1973), .B(n1975), .CI(n1971), .CO(n1955), .S(n1956) );
  FA_X1 U1348 ( .A(n2493), .B(n2557), .CI(n2525), .CO(n1957), .S(n1958) );
  FA_X1 U1349 ( .A(n2429), .B(n2589), .CI(n2461), .CO(n1959), .S(n1960) );
  FA_X1 U1350 ( .A(n2397), .B(n2621), .CI(n2365), .CO(n1961), .S(n1962) );
  FA_X1 U1351 ( .A(n1979), .B(n1968), .CI(n1966), .CO(n1963), .S(n1964) );
  FA_X1 U1352 ( .A(n1981), .B(n1974), .CI(n1970), .CO(n1965), .S(n1966) );
  FA_X1 U1353 ( .A(n1983), .B(n1985), .CI(n1972), .CO(n1967), .S(n1968) );
  FA_X1 U1354 ( .A(n1976), .B(n2494), .CI(n1987), .CO(n1969), .S(n1970) );
  FA_X1 U1355 ( .A(n2558), .B(n2430), .CI(n2462), .CO(n1971), .S(n1972) );
  FA_X1 U1356 ( .A(n2622), .B(n2526), .CI(n2590), .CO(n1973), .S(n1974) );
  HA_X1 U1357 ( .A(n2398), .B(n2069), .CO(n1975), .S(n1976) );
  FA_X1 U1358 ( .A(n1991), .B(n1982), .CI(n1980), .CO(n1977), .S(n1978) );
  FA_X1 U1359 ( .A(n1984), .B(n1988), .CI(n1993), .CO(n1979), .S(n1980) );
  FA_X1 U1360 ( .A(n1995), .B(n1997), .CI(n1986), .CO(n1981), .S(n1982) );
  FA_X1 U1361 ( .A(n2527), .B(n2559), .CI(n1999), .CO(n1983), .S(n1984) );
  FA_X1 U1362 ( .A(n2463), .B(n2591), .CI(n2495), .CO(n1985), .S(n1986) );
  FA_X1 U1363 ( .A(n2431), .B(n2623), .CI(n2399), .CO(n1987), .S(n1988) );
  FA_X1 U1364 ( .A(n2003), .B(n1994), .CI(n1992), .CO(n1989), .S(n1990) );
  FA_X1 U1365 ( .A(n1998), .B(n1996), .CI(n2005), .CO(n1991), .S(n1992) );
  FA_X1 U1366 ( .A(n2009), .B(n2000), .CI(n2007), .CO(n1993), .S(n1994) );
  FA_X1 U1367 ( .A(n2464), .B(n2560), .CI(n2496), .CO(n1995), .S(n1996) );
  FA_X1 U1368 ( .A(n2624), .B(n2528), .CI(n2592), .CO(n1997), .S(n1998) );
  HA_X1 U1369 ( .A(n2432), .B(n2070), .CO(n1999), .S(n2000) );
  FA_X1 U1370 ( .A(n2006), .B(n2013), .CI(n2004), .CO(n2001), .S(n2002) );
  FA_X1 U1371 ( .A(n2010), .B(n2008), .CI(n2015), .CO(n2003), .S(n2004) );
  FA_X1 U1372 ( .A(n2019), .B(n2561), .CI(n2017), .CO(n2005), .S(n2006) );
  FA_X1 U1373 ( .A(n2497), .B(n2593), .CI(n2529), .CO(n2007), .S(n2008) );
  FA_X1 U1374 ( .A(n2465), .B(n2625), .CI(n2433), .CO(n2009), .S(n2010) );
  FA_X1 U1375 ( .A(n2023), .B(n2016), .CI(n2014), .CO(n2011), .S(n2012) );
  FA_X1 U1376 ( .A(n2025), .B(n2027), .CI(n2018), .CO(n2013), .S(n2014) );
  FA_X1 U1377 ( .A(n2498), .B(n2530), .CI(n2020), .CO(n2015), .S(n2016) );
  FA_X1 U1378 ( .A(n2626), .B(n2562), .CI(n2594), .CO(n2017), .S(n2018) );
  HA_X1 U1379 ( .A(n2466), .B(n2071), .CO(n2019), .S(n2020) );
  FA_X1 U1380 ( .A(n2031), .B(n2028), .CI(n2024), .CO(n2021), .S(n2022) );
  FA_X1 U1381 ( .A(n2033), .B(n2035), .CI(n2026), .CO(n2023), .S(n2024) );
  FA_X1 U1382 ( .A(n2531), .B(n2595), .CI(n2563), .CO(n2025), .S(n2026) );
  FA_X1 U1383 ( .A(n2499), .B(n2627), .CI(n2467), .CO(n2027), .S(n2028) );
  FA_X1 U1384 ( .A(n2034), .B(n2039), .CI(n2032), .CO(n2029), .S(n2030) );
  FA_X1 U1385 ( .A(n2036), .B(n2628), .CI(n2041), .CO(n2031), .S(n2032) );
  FA_X1 U1386 ( .A(n2532), .B(n2564), .CI(n2596), .CO(n2033), .S(n2034) );
  HA_X1 U1387 ( .A(n2500), .B(n2072), .CO(n2035), .S(n2036) );
  FA_X1 U1388 ( .A(n2042), .B(n2045), .CI(n2040), .CO(n2037), .S(n2038) );
  FA_X1 U1389 ( .A(n2565), .B(n2597), .CI(n2047), .CO(n2039), .S(n2040) );
  FA_X1 U1390 ( .A(n2533), .B(n2629), .CI(n2501), .CO(n2041), .S(n2042) );
  FA_X1 U1391 ( .A(n2051), .B(n2048), .CI(n2046), .CO(n2043), .S(n2044) );
  FA_X1 U1392 ( .A(n2566), .B(n2630), .CI(n2598), .CO(n2045), .S(n2046) );
  HA_X1 U1393 ( .A(n2534), .B(n2073), .CO(n2047), .S(n2048) );
  FA_X1 U1394 ( .A(n2055), .B(n2599), .CI(n2052), .CO(n2049), .S(n2050) );
  FA_X1 U1395 ( .A(n2567), .B(n2631), .CI(n2535), .CO(n2051), .S(n2052) );
  FA_X1 U1396 ( .A(n2600), .B(n2632), .CI(n2056), .CO(n2053), .S(n2054) );
  HA_X1 U1397 ( .A(n2568), .B(n2074), .CO(n2055), .S(n2056) );
  FA_X1 U1398 ( .A(n2601), .B(n2633), .CI(n2569), .CO(n2057), .S(n2058) );
  HA_X1 U1399 ( .A(n2634), .B(n2602), .CO(n2059), .S(n2060) );
  NOR2_X4 U1400 ( .A1(n2637), .A2(n3455), .ZN(n2077) );
  NOR2_X4 U1401 ( .A1(n2638), .A2(n3455), .ZN(n1044) );
  NOR2_X4 U1402 ( .A1(n2639), .A2(n3455), .ZN(n2078) );
  NOR2_X4 U1403 ( .A1(n2640), .A2(n3455), .ZN(n1054) );
  NOR2_X4 U1404 ( .A1(n2641), .A2(n3455), .ZN(n2079) );
  NOR2_X4 U1405 ( .A1(n2642), .A2(n3455), .ZN(n1068) );
  NOR2_X4 U1406 ( .A1(n2643), .A2(n3455), .ZN(n2080) );
  NOR2_X4 U1407 ( .A1(n2644), .A2(n3455), .ZN(n1086) );
  NOR2_X4 U1408 ( .A1(n2645), .A2(n3455), .ZN(n2081) );
  NOR2_X4 U1409 ( .A1(n2646), .A2(n3455), .ZN(n1108) );
  NOR2_X4 U1410 ( .A1(n2647), .A2(n3455), .ZN(n2082) );
  NOR2_X4 U1411 ( .A1(n2648), .A2(n3455), .ZN(n1134) );
  NOR2_X4 U1412 ( .A1(n2649), .A2(n3455), .ZN(n2083) );
  NOR2_X4 U1413 ( .A1(n2650), .A2(n3455), .ZN(n1164) );
  NOR2_X4 U1414 ( .A1(n2651), .A2(n3455), .ZN(n2084) );
  NOR2_X4 U1415 ( .A1(n2652), .A2(n3455), .ZN(n1198) );
  NOR2_X4 U1416 ( .A1(n2653), .A2(n3455), .ZN(n2085) );
  NOR2_X4 U1417 ( .A1(n2654), .A2(n3455), .ZN(n1236) );
  NOR2_X4 U1418 ( .A1(n2655), .A2(n3455), .ZN(n2086) );
  NOR2_X4 U1419 ( .A1(n2656), .A2(n3455), .ZN(n1278) );
  NOR2_X4 U1420 ( .A1(n2657), .A2(n3455), .ZN(n2087) );
  NOR2_X4 U1421 ( .A1(n2658), .A2(n3455), .ZN(n1324) );
  NOR2_X4 U1422 ( .A1(n2659), .A2(n3455), .ZN(n2088) );
  NOR2_X4 U1423 ( .A1(n2660), .A2(n3455), .ZN(n1374) );
  NOR2_X4 U1424 ( .A1(n2661), .A2(n3455), .ZN(n2089) );
  NOR2_X4 U1426 ( .A1(n2663), .A2(n3455), .ZN(n2090) );
  NOR2_X4 U1427 ( .A1(n2664), .A2(n3455), .ZN(n1486) );
  NOR2_X4 U1428 ( .A1(n2665), .A2(n3455), .ZN(n2091) );
  NOR2_X4 U1429 ( .A1(n2666), .A2(n3455), .ZN(n2092) );
  NOR2_X4 U1430 ( .A1(n2667), .A2(n3455), .ZN(n1548) );
  OAI22_X2 U1462 ( .A1(n464), .A2(n3455), .B1(n2700), .B2(n3526), .ZN(n2061)
         );
  OAI22_X2 U1463 ( .A1(n3525), .A2(n2668), .B1(n3526), .B2(n3455), .ZN(n2095)
         );
  OAI22_X2 U1464 ( .A1(n3525), .A2(n2669), .B1(n2668), .B2(n3526), .ZN(n2096)
         );
  OAI22_X2 U1465 ( .A1(n3525), .A2(n2670), .B1(n2669), .B2(n3526), .ZN(n2097)
         );
  OAI22_X2 U1466 ( .A1(n3525), .A2(n2671), .B1(n2670), .B2(n3526), .ZN(n2098)
         );
  OAI22_X2 U1467 ( .A1(n3525), .A2(n2672), .B1(n2671), .B2(n3526), .ZN(n2099)
         );
  OAI22_X2 U1468 ( .A1(n3525), .A2(n2673), .B1(n2672), .B2(n3526), .ZN(n2100)
         );
  OAI22_X2 U1469 ( .A1(n3525), .A2(n2674), .B1(n2673), .B2(n3526), .ZN(n2101)
         );
  OAI22_X2 U1470 ( .A1(n3525), .A2(n2675), .B1(n2674), .B2(n3526), .ZN(n2102)
         );
  OAI22_X2 U1471 ( .A1(n464), .A2(n2676), .B1(n2675), .B2(n3526), .ZN(n2103)
         );
  OAI22_X2 U1472 ( .A1(n464), .A2(n2677), .B1(n2676), .B2(n3526), .ZN(n2104)
         );
  OAI22_X2 U1473 ( .A1(n464), .A2(n2678), .B1(n2677), .B2(n3526), .ZN(n2105)
         );
  OAI22_X2 U1474 ( .A1(n464), .A2(n2679), .B1(n2678), .B2(n3526), .ZN(n2106)
         );
  OAI22_X2 U1475 ( .A1(n464), .A2(n2680), .B1(n2679), .B2(n3526), .ZN(n2107)
         );
  OAI22_X2 U1476 ( .A1(n464), .A2(n2681), .B1(n2680), .B2(n3526), .ZN(n2108)
         );
  OAI22_X2 U1477 ( .A1(n464), .A2(n2682), .B1(n2681), .B2(n3526), .ZN(n2109)
         );
  OAI22_X2 U1478 ( .A1(n464), .A2(n2683), .B1(n2682), .B2(n3526), .ZN(n2110)
         );
  OAI22_X2 U1479 ( .A1(n464), .A2(n2684), .B1(n2683), .B2(n3526), .ZN(n2111)
         );
  OAI22_X2 U1480 ( .A1(n464), .A2(n2685), .B1(n2684), .B2(n3526), .ZN(n2112)
         );
  OAI22_X2 U1481 ( .A1(n464), .A2(n2686), .B1(n2685), .B2(n3526), .ZN(n2113)
         );
  OAI22_X2 U1482 ( .A1(n464), .A2(n2687), .B1(n2686), .B2(n3526), .ZN(n2114)
         );
  OAI22_X2 U1483 ( .A1(n464), .A2(n2688), .B1(n2687), .B2(n3526), .ZN(n2115)
         );
  OAI22_X2 U1484 ( .A1(n464), .A2(n2689), .B1(n2688), .B2(n3526), .ZN(n2116)
         );
  OAI22_X2 U1485 ( .A1(n464), .A2(n2690), .B1(n2689), .B2(n3526), .ZN(n2117)
         );
  OAI22_X2 U1487 ( .A1(n464), .A2(n2692), .B1(n2691), .B2(n3526), .ZN(n2119)
         );
  OAI22_X2 U1489 ( .A1(n464), .A2(n2694), .B1(n2693), .B2(n3526), .ZN(n2121)
         );
  OAI22_X2 U1490 ( .A1(n464), .A2(n2695), .B1(n2694), .B2(n3526), .ZN(n2122)
         );
  OAI22_X2 U1493 ( .A1(n464), .A2(n2698), .B1(n2697), .B2(n3526), .ZN(n2125)
         );
  OAI22_X2 U1528 ( .A1(n3476), .A2(n2701), .B1(n3557), .B2(n3278), .ZN(n2129)
         );
  OAI22_X2 U1530 ( .A1(n3476), .A2(n2703), .B1(n2702), .B2(n3557), .ZN(n2131)
         );
  OAI22_X2 U1531 ( .A1(n3476), .A2(n2704), .B1(n2703), .B2(n3557), .ZN(n2132)
         );
  OAI22_X2 U1533 ( .A1(n3476), .A2(n2706), .B1(n2705), .B2(n3557), .ZN(n2134)
         );
  OAI22_X2 U1539 ( .A1(n3476), .A2(n2712), .B1(n2711), .B2(n3557), .ZN(n2140)
         );
  OAI22_X2 U1541 ( .A1(n461), .A2(n2714), .B1(n2713), .B2(n3557), .ZN(n2142)
         );
  OAI22_X2 U1543 ( .A1(n3476), .A2(n2716), .B1(n2715), .B2(n3557), .ZN(n2144)
         );
  OAI22_X2 U1544 ( .A1(n3476), .A2(n2717), .B1(n2716), .B2(n3557), .ZN(n2145)
         );
  OAI22_X2 U1545 ( .A1(n3476), .A2(n2718), .B1(n2717), .B2(n3557), .ZN(n2146)
         );
  OAI22_X2 U1546 ( .A1(n3476), .A2(n2719), .B1(n2718), .B2(n3557), .ZN(n2147)
         );
  OAI22_X2 U1548 ( .A1(n3476), .A2(n2721), .B1(n2720), .B2(n3557), .ZN(n2149)
         );
  OAI22_X2 U1593 ( .A1(n3506), .A2(n2734), .B1(n408), .B2(n3279), .ZN(n2163)
         );
  OAI22_X2 U1594 ( .A1(n3506), .A2(n2735), .B1(n2734), .B2(n408), .ZN(n2164)
         );
  OAI22_X2 U1595 ( .A1(n3506), .A2(n2736), .B1(n2735), .B2(n408), .ZN(n2165)
         );
  OAI22_X2 U1596 ( .A1(n3506), .A2(n2737), .B1(n2736), .B2(n408), .ZN(n2166)
         );
  OAI22_X2 U1597 ( .A1(n3506), .A2(n2738), .B1(n2737), .B2(n408), .ZN(n2167)
         );
  OAI22_X2 U1599 ( .A1(n3506), .A2(n2740), .B1(n2739), .B2(n408), .ZN(n2169)
         );
  OAI22_X2 U1600 ( .A1(n3506), .A2(n2741), .B1(n2740), .B2(n408), .ZN(n2170)
         );
  OAI22_X2 U1601 ( .A1(n3506), .A2(n2742), .B1(n2741), .B2(n408), .ZN(n2171)
         );
  OAI22_X2 U1602 ( .A1(n3506), .A2(n2743), .B1(n2742), .B2(n408), .ZN(n2172)
         );
  OAI22_X2 U1603 ( .A1(n3506), .A2(n2744), .B1(n2743), .B2(n408), .ZN(n2173)
         );
  OAI22_X2 U1606 ( .A1(n3506), .A2(n2747), .B1(n2746), .B2(n408), .ZN(n2176)
         );
  OAI22_X2 U1608 ( .A1(n3506), .A2(n2749), .B1(n2748), .B2(n408), .ZN(n2178)
         );
  OAI22_X2 U1609 ( .A1(n3506), .A2(n2750), .B1(n2749), .B2(n408), .ZN(n2179)
         );
  OAI22_X2 U1610 ( .A1(n3506), .A2(n2751), .B1(n2750), .B2(n408), .ZN(n2180)
         );
  OAI22_X2 U1611 ( .A1(n3506), .A2(n2752), .B1(n2751), .B2(n408), .ZN(n2181)
         );
  OAI22_X2 U1616 ( .A1(n3506), .A2(n2757), .B1(n2756), .B2(n408), .ZN(n2186)
         );
  OAI22_X2 U1624 ( .A1(n3506), .A2(n2765), .B1(n2764), .B2(n408), .ZN(n2194)
         );
  OAI22_X2 U1722 ( .A1(n3671), .A2(n3281), .B1(n2832), .B2(n402), .ZN(n2065)
         );
  OAI22_X2 U1723 ( .A1(n3671), .A2(n2800), .B1(n402), .B2(n3281), .ZN(n2231)
         );
  OAI22_X2 U1724 ( .A1(n3671), .A2(n2801), .B1(n2800), .B2(n402), .ZN(n2232)
         );
  OAI22_X2 U1725 ( .A1(n3671), .A2(n2802), .B1(n2801), .B2(n402), .ZN(n2233)
         );
  OAI22_X2 U1726 ( .A1(n3671), .A2(n2803), .B1(n2802), .B2(n402), .ZN(n2234)
         );
  OAI22_X2 U1727 ( .A1(n3671), .A2(n2804), .B1(n2803), .B2(n402), .ZN(n2235)
         );
  OAI22_X2 U1729 ( .A1(n3671), .A2(n2806), .B1(n2805), .B2(n402), .ZN(n2237)
         );
  OAI22_X2 U1730 ( .A1(n452), .A2(n2807), .B1(n2806), .B2(n402), .ZN(n2238) );
  OAI22_X2 U1731 ( .A1(n3671), .A2(n2808), .B1(n2807), .B2(n402), .ZN(n2239)
         );
  OAI22_X2 U1732 ( .A1(n3671), .A2(n2809), .B1(n2808), .B2(n402), .ZN(n2240)
         );
  OAI22_X2 U1733 ( .A1(n452), .A2(n2810), .B1(n2809), .B2(n402), .ZN(n2241) );
  OAI22_X2 U1736 ( .A1(n3671), .A2(n2813), .B1(n2812), .B2(n402), .ZN(n2244)
         );
  OAI22_X2 U1737 ( .A1(n3671), .A2(n2814), .B1(n2813), .B2(n402), .ZN(n2245)
         );
  OAI22_X2 U1739 ( .A1(n3671), .A2(n2816), .B1(n2815), .B2(n402), .ZN(n2247)
         );
  OAI22_X2 U1750 ( .A1(n3671), .A2(n2827), .B1(n2826), .B2(n402), .ZN(n2258)
         );
  OAI22_X2 U1754 ( .A1(n3671), .A2(n2831), .B1(n2830), .B2(n402), .ZN(n2262)
         );
  OAI22_X2 U1787 ( .A1(n449), .A2(n3282), .B1(n2865), .B2(n399), .ZN(n2066) );
  OAI22_X2 U1788 ( .A1(n449), .A2(n2833), .B1(n399), .B2(n3282), .ZN(n2265) );
  OAI22_X2 U1789 ( .A1(n449), .A2(n2834), .B1(n2833), .B2(n399), .ZN(n2266) );
  OAI22_X2 U1790 ( .A1(n449), .A2(n2835), .B1(n2834), .B2(n399), .ZN(n2267) );
  OAI22_X2 U1791 ( .A1(n449), .A2(n2836), .B1(n2835), .B2(n399), .ZN(n2268) );
  OAI22_X2 U1792 ( .A1(n449), .A2(n2837), .B1(n2836), .B2(n399), .ZN(n2269) );
  OAI22_X2 U1793 ( .A1(n449), .A2(n2838), .B1(n2837), .B2(n399), .ZN(n2270) );
  OAI22_X2 U1795 ( .A1(n449), .A2(n2840), .B1(n2839), .B2(n399), .ZN(n2272) );
  OAI22_X2 U1796 ( .A1(n449), .A2(n2841), .B1(n2840), .B2(n399), .ZN(n2273) );
  OAI22_X2 U1797 ( .A1(n449), .A2(n2842), .B1(n2841), .B2(n399), .ZN(n2274) );
  OAI22_X2 U1798 ( .A1(n449), .A2(n2843), .B1(n2842), .B2(n399), .ZN(n2275) );
  OAI22_X2 U1799 ( .A1(n449), .A2(n2844), .B1(n2843), .B2(n399), .ZN(n2276) );
  OAI22_X2 U1800 ( .A1(n449), .A2(n2845), .B1(n2844), .B2(n399), .ZN(n2277) );
  OAI22_X2 U1802 ( .A1(n449), .A2(n2847), .B1(n2846), .B2(n399), .ZN(n2279) );
  OAI22_X2 U1804 ( .A1(n449), .A2(n2849), .B1(n2848), .B2(n399), .ZN(n2281) );
  OAI22_X2 U1805 ( .A1(n449), .A2(n2850), .B1(n2849), .B2(n399), .ZN(n2282) );
  OAI22_X2 U1806 ( .A1(n449), .A2(n2851), .B1(n2850), .B2(n399), .ZN(n2283) );
  OAI22_X2 U1807 ( .A1(n449), .A2(n2852), .B1(n2851), .B2(n399), .ZN(n2284) );
  OAI22_X2 U1808 ( .A1(n449), .A2(n2853), .B1(n2852), .B2(n399), .ZN(n2285) );
  OAI22_X2 U1809 ( .A1(n449), .A2(n2854), .B1(n2853), .B2(n399), .ZN(n2286) );
  OAI22_X2 U1810 ( .A1(n449), .A2(n2855), .B1(n2854), .B2(n399), .ZN(n2287) );
  OAI22_X2 U1812 ( .A1(n449), .A2(n2857), .B1(n2856), .B2(n399), .ZN(n2289) );
  OAI22_X2 U1813 ( .A1(n449), .A2(n2858), .B1(n2857), .B2(n399), .ZN(n2290) );
  OAI22_X2 U1814 ( .A1(n449), .A2(n2859), .B1(n2858), .B2(n399), .ZN(n2291) );
  OAI22_X2 U1816 ( .A1(n449), .A2(n2861), .B1(n2860), .B2(n399), .ZN(n2293) );
  OAI22_X2 U1817 ( .A1(n449), .A2(n2862), .B1(n2861), .B2(n399), .ZN(n2294) );
  OAI22_X2 U1819 ( .A1(n449), .A2(n2864), .B1(n2863), .B2(n399), .ZN(n2296) );
  OAI22_X2 U1853 ( .A1(n3666), .A2(n2866), .B1(n396), .B2(n3283), .ZN(n2299)
         );
  OAI22_X2 U1854 ( .A1(n3666), .A2(n2867), .B1(n2866), .B2(n396), .ZN(n2300)
         );
  OAI22_X2 U1855 ( .A1(n3666), .A2(n2868), .B1(n2867), .B2(n396), .ZN(n2301)
         );
  OAI22_X2 U1856 ( .A1(n3666), .A2(n2869), .B1(n2868), .B2(n396), .ZN(n2302)
         );
  OAI22_X2 U1857 ( .A1(n3666), .A2(n2870), .B1(n2869), .B2(n396), .ZN(n2303)
         );
  OAI22_X2 U1858 ( .A1(n3666), .A2(n2871), .B1(n2870), .B2(n396), .ZN(n2304)
         );
  OAI22_X2 U1859 ( .A1(n3666), .A2(n2872), .B1(n2871), .B2(n396), .ZN(n2305)
         );
  OAI22_X2 U1860 ( .A1(n3666), .A2(n2873), .B1(n2872), .B2(n396), .ZN(n2306)
         );
  OAI22_X2 U1861 ( .A1(n3666), .A2(n2874), .B1(n2873), .B2(n396), .ZN(n2307)
         );
  OAI22_X2 U1862 ( .A1(n3666), .A2(n2875), .B1(n2874), .B2(n396), .ZN(n2308)
         );
  OAI22_X2 U1863 ( .A1(n3666), .A2(n2876), .B1(n2875), .B2(n396), .ZN(n2309)
         );
  OAI22_X2 U1865 ( .A1(n3666), .A2(n2878), .B1(n2877), .B2(n396), .ZN(n2311)
         );
  OAI22_X2 U1873 ( .A1(n3666), .A2(n2886), .B1(n2885), .B2(n396), .ZN(n2319)
         );
  OAI22_X2 U1876 ( .A1(n3666), .A2(n2889), .B1(n2888), .B2(n396), .ZN(n2322)
         );
  OAI22_X2 U1877 ( .A1(n3666), .A2(n2890), .B1(n2889), .B2(n396), .ZN(n2323)
         );
  OAI22_X2 U1878 ( .A1(n3666), .A2(n2891), .B1(n2890), .B2(n396), .ZN(n2324)
         );
  OAI22_X2 U1879 ( .A1(n3666), .A2(n2892), .B1(n2891), .B2(n396), .ZN(n2325)
         );
  OAI22_X2 U1880 ( .A1(n3666), .A2(n2893), .B1(n2892), .B2(n396), .ZN(n2326)
         );
  OAI22_X2 U1881 ( .A1(n3666), .A2(n2894), .B1(n2893), .B2(n396), .ZN(n2327)
         );
  OAI22_X2 U1882 ( .A1(n3666), .A2(n2895), .B1(n2894), .B2(n396), .ZN(n2328)
         );
  OAI22_X2 U1884 ( .A1(n3666), .A2(n2897), .B1(n2896), .B2(n396), .ZN(n2330)
         );
  OAI22_X2 U1918 ( .A1(n3650), .A2(n2899), .B1(n3556), .B2(n3284), .ZN(n2333)
         );
  OAI22_X2 U1920 ( .A1(n3650), .A2(n2901), .B1(n2900), .B2(n3556), .ZN(n2335)
         );
  OAI22_X2 U1922 ( .A1(n3650), .A2(n2903), .B1(n2902), .B2(n3556), .ZN(n2337)
         );
  OAI22_X2 U1923 ( .A1(n3650), .A2(n2904), .B1(n2903), .B2(n3556), .ZN(n2338)
         );
  OAI22_X2 U1926 ( .A1(n3650), .A2(n2907), .B1(n2906), .B2(n3556), .ZN(n2341)
         );
  OAI22_X2 U1927 ( .A1(n3649), .A2(n2908), .B1(n2907), .B2(n3556), .ZN(n2342)
         );
  OAI22_X2 U1928 ( .A1(n3650), .A2(n2909), .B1(n2908), .B2(n3556), .ZN(n2343)
         );
  OAI22_X2 U1930 ( .A1(n3650), .A2(n2911), .B1(n2910), .B2(n3556), .ZN(n2345)
         );
  OAI22_X2 U1933 ( .A1(n3649), .A2(n2914), .B1(n2913), .B2(n3556), .ZN(n2348)
         );
  OAI22_X2 U1935 ( .A1(n3650), .A2(n2916), .B1(n2915), .B2(n3556), .ZN(n2350)
         );
  OAI22_X2 U1937 ( .A1(n3650), .A2(n2918), .B1(n2917), .B2(n3556), .ZN(n2352)
         );
  OAI22_X2 U1943 ( .A1(n3650), .A2(n2924), .B1(n2923), .B2(n3556), .ZN(n2358)
         );
  OAI22_X2 U1982 ( .A1(n440), .A2(n3285), .B1(n2964), .B2(n390), .ZN(n2069) );
  OAI22_X2 U1983 ( .A1(n3535), .A2(n2932), .B1(n390), .B2(n3285), .ZN(n2367)
         );
  OAI22_X2 U1984 ( .A1(n3535), .A2(n2933), .B1(n2932), .B2(n390), .ZN(n2368)
         );
  OAI22_X2 U1985 ( .A1(n3535), .A2(n2934), .B1(n2933), .B2(n390), .ZN(n2369)
         );
  OAI22_X2 U1986 ( .A1(n3535), .A2(n2935), .B1(n2934), .B2(n390), .ZN(n2370)
         );
  OAI22_X2 U1987 ( .A1(n440), .A2(n2936), .B1(n2935), .B2(n390), .ZN(n2371) );
  OAI22_X2 U1988 ( .A1(n3535), .A2(n2937), .B1(n2936), .B2(n390), .ZN(n2372)
         );
  OAI22_X2 U1989 ( .A1(n3535), .A2(n2938), .B1(n2937), .B2(n390), .ZN(n2373)
         );
  OAI22_X2 U1990 ( .A1(n3535), .A2(n2939), .B1(n2938), .B2(n390), .ZN(n2374)
         );
  OAI22_X2 U1992 ( .A1(n3535), .A2(n2941), .B1(n2940), .B2(n390), .ZN(n2376)
         );
  OAI22_X2 U1993 ( .A1(n3535), .A2(n2942), .B1(n2941), .B2(n390), .ZN(n2377)
         );
  OAI22_X2 U1994 ( .A1(n440), .A2(n2943), .B1(n2942), .B2(n390), .ZN(n2378) );
  OAI22_X2 U1995 ( .A1(n440), .A2(n2944), .B1(n2943), .B2(n390), .ZN(n2379) );
  OAI22_X2 U1996 ( .A1(n440), .A2(n2945), .B1(n2944), .B2(n390), .ZN(n2380) );
  OAI22_X2 U1997 ( .A1(n440), .A2(n2946), .B1(n2945), .B2(n390), .ZN(n2381) );
  OAI22_X2 U1998 ( .A1(n440), .A2(n2947), .B1(n2946), .B2(n390), .ZN(n2382) );
  OAI22_X2 U1999 ( .A1(n3535), .A2(n2948), .B1(n2947), .B2(n390), .ZN(n2383)
         );
  OAI22_X2 U2000 ( .A1(n440), .A2(n2949), .B1(n2948), .B2(n390), .ZN(n2384) );
  OAI22_X2 U2001 ( .A1(n3535), .A2(n2950), .B1(n2949), .B2(n390), .ZN(n2385)
         );
  OAI22_X2 U2002 ( .A1(n440), .A2(n2951), .B1(n2950), .B2(n390), .ZN(n2386) );
  OAI22_X2 U2003 ( .A1(n3535), .A2(n2952), .B1(n2951), .B2(n390), .ZN(n2387)
         );
  OAI22_X2 U2004 ( .A1(n440), .A2(n2953), .B1(n2952), .B2(n390), .ZN(n2388) );
  OAI22_X2 U2005 ( .A1(n440), .A2(n2954), .B1(n2953), .B2(n390), .ZN(n2389) );
  OAI22_X2 U2006 ( .A1(n440), .A2(n2955), .B1(n2954), .B2(n390), .ZN(n2390) );
  OAI22_X2 U2007 ( .A1(n440), .A2(n2956), .B1(n2955), .B2(n390), .ZN(n2391) );
  OAI22_X2 U2008 ( .A1(n3535), .A2(n2957), .B1(n2956), .B2(n390), .ZN(n2392)
         );
  OAI22_X2 U2009 ( .A1(n3535), .A2(n2958), .B1(n2957), .B2(n390), .ZN(n2393)
         );
  OAI22_X2 U2010 ( .A1(n440), .A2(n2959), .B1(n2958), .B2(n390), .ZN(n2394) );
  OAI22_X2 U2011 ( .A1(n3535), .A2(n2960), .B1(n2959), .B2(n390), .ZN(n2395)
         );
  OAI22_X2 U2012 ( .A1(n440), .A2(n2961), .B1(n2960), .B2(n390), .ZN(n2396) );
  OAI22_X2 U2013 ( .A1(n3535), .A2(n2962), .B1(n2961), .B2(n390), .ZN(n2397)
         );
  OAI22_X2 U2014 ( .A1(n440), .A2(n2963), .B1(n2962), .B2(n390), .ZN(n2398) );
  OAI22_X2 U2047 ( .A1(n3436), .A2(n3286), .B1(n2997), .B2(n387), .ZN(n2070)
         );
  OAI22_X2 U2048 ( .A1(n3436), .A2(n2965), .B1(n387), .B2(n3286), .ZN(n2401)
         );
  OAI22_X2 U2049 ( .A1(n3436), .A2(n2966), .B1(n2965), .B2(n387), .ZN(n2402)
         );
  OAI22_X2 U2050 ( .A1(n3435), .A2(n2967), .B1(n2966), .B2(n387), .ZN(n2403)
         );
  OAI22_X2 U2051 ( .A1(n3436), .A2(n2968), .B1(n2967), .B2(n387), .ZN(n2404)
         );
  OAI22_X2 U2052 ( .A1(n3435), .A2(n2969), .B1(n2968), .B2(n387), .ZN(n2405)
         );
  OAI22_X2 U2055 ( .A1(n3435), .A2(n2972), .B1(n2971), .B2(n387), .ZN(n2408)
         );
  OAI22_X2 U2056 ( .A1(n3436), .A2(n2973), .B1(n2972), .B2(n387), .ZN(n2409)
         );
  OAI22_X2 U2057 ( .A1(n3436), .A2(n2974), .B1(n2973), .B2(n387), .ZN(n2410)
         );
  OAI22_X2 U2058 ( .A1(n3435), .A2(n2975), .B1(n2974), .B2(n387), .ZN(n2411)
         );
  OAI22_X2 U2060 ( .A1(n3435), .A2(n2977), .B1(n2976), .B2(n387), .ZN(n2413)
         );
  OAI22_X2 U2061 ( .A1(n3436), .A2(n2978), .B1(n2977), .B2(n387), .ZN(n2414)
         );
  OAI22_X2 U2063 ( .A1(n3435), .A2(n2980), .B1(n2979), .B2(n387), .ZN(n2416)
         );
  OAI22_X2 U2064 ( .A1(n3435), .A2(n2981), .B1(n2980), .B2(n387), .ZN(n2417)
         );
  OAI22_X2 U2065 ( .A1(n3435), .A2(n2982), .B1(n2981), .B2(n387), .ZN(n2418)
         );
  OAI22_X2 U2068 ( .A1(n437), .A2(n2985), .B1(n2984), .B2(n387), .ZN(n2421) );
  OAI22_X2 U2069 ( .A1(n3435), .A2(n2986), .B1(n2985), .B2(n387), .ZN(n2422)
         );
  OAI22_X2 U2070 ( .A1(n3435), .A2(n2987), .B1(n2986), .B2(n387), .ZN(n2423)
         );
  OAI22_X2 U2071 ( .A1(n3436), .A2(n2988), .B1(n2987), .B2(n387), .ZN(n2424)
         );
  OAI22_X2 U2073 ( .A1(n3435), .A2(n2990), .B1(n2989), .B2(n387), .ZN(n2426)
         );
  OAI22_X2 U2074 ( .A1(n3436), .A2(n2991), .B1(n2990), .B2(n387), .ZN(n2427)
         );
  OAI22_X2 U2075 ( .A1(n3436), .A2(n2992), .B1(n2991), .B2(n387), .ZN(n2428)
         );
  OAI22_X2 U2076 ( .A1(n3436), .A2(n2993), .B1(n2992), .B2(n387), .ZN(n2429)
         );
  OAI22_X2 U2077 ( .A1(n3436), .A2(n2994), .B1(n2993), .B2(n387), .ZN(n2430)
         );
  OAI22_X2 U2078 ( .A1(n3435), .A2(n2995), .B1(n2994), .B2(n387), .ZN(n2431)
         );
  OAI22_X2 U2079 ( .A1(n3436), .A2(n2996), .B1(n2995), .B2(n387), .ZN(n2432)
         );
  OAI22_X2 U2311 ( .A1(n3537), .A2(n3100), .B1(n3099), .B2(n375), .ZN(n2540)
         );
  OAI22_X2 U2437 ( .A1(n419), .A2(n3292), .B1(n3195), .B2(n369), .ZN(n2076) );
  OAI22_X2 U2438 ( .A1(n419), .A2(n3163), .B1(n3292), .B2(n369), .ZN(n2605) );
  OAI22_X2 U2439 ( .A1(n419), .A2(n3164), .B1(n3163), .B2(n369), .ZN(n2606) );
  OAI22_X2 U2441 ( .A1(n419), .A2(n3166), .B1(n3165), .B2(n369), .ZN(n2608) );
  OAI22_X2 U2442 ( .A1(n419), .A2(n3167), .B1(n3166), .B2(n369), .ZN(n2609) );
  OAI22_X2 U2443 ( .A1(n419), .A2(n3168), .B1(n3167), .B2(n369), .ZN(n2610) );
  OAI22_X2 U2444 ( .A1(n419), .A2(n3169), .B1(n3168), .B2(n369), .ZN(n2611) );
  OAI22_X2 U2445 ( .A1(n419), .A2(n3170), .B1(n3169), .B2(n369), .ZN(n2612) );
  OAI22_X2 U2446 ( .A1(n419), .A2(n3171), .B1(n3170), .B2(n369), .ZN(n2613) );
  OAI22_X2 U2447 ( .A1(n419), .A2(n3172), .B1(n3171), .B2(n369), .ZN(n2614) );
  OAI22_X2 U2448 ( .A1(n419), .A2(n3173), .B1(n3172), .B2(n369), .ZN(n2615) );
  OAI22_X2 U2449 ( .A1(n419), .A2(n3174), .B1(n3173), .B2(n369), .ZN(n2616) );
  OAI22_X2 U2450 ( .A1(n419), .A2(n3175), .B1(n3174), .B2(n369), .ZN(n2617) );
  OAI22_X2 U2451 ( .A1(n419), .A2(n3176), .B1(n3175), .B2(n369), .ZN(n2618) );
  OAI22_X2 U2452 ( .A1(n419), .A2(n3177), .B1(n3176), .B2(n369), .ZN(n2619) );
  OAI22_X2 U2453 ( .A1(n419), .A2(n3178), .B1(n3177), .B2(n369), .ZN(n2620) );
  OAI22_X2 U2454 ( .A1(n419), .A2(n3179), .B1(n3178), .B2(n369), .ZN(n2621) );
  OAI22_X2 U2455 ( .A1(n419), .A2(n3180), .B1(n3179), .B2(n369), .ZN(n2622) );
  OAI22_X2 U2456 ( .A1(n419), .A2(n3181), .B1(n3180), .B2(n369), .ZN(n2623) );
  OAI22_X2 U2457 ( .A1(n419), .A2(n3182), .B1(n3181), .B2(n369), .ZN(n2624) );
  OAI22_X2 U2458 ( .A1(n419), .A2(n3183), .B1(n3182), .B2(n369), .ZN(n2625) );
  OAI22_X2 U2459 ( .A1(n419), .A2(n3184), .B1(n3183), .B2(n369), .ZN(n2626) );
  OAI22_X2 U2460 ( .A1(n419), .A2(n3185), .B1(n3184), .B2(n369), .ZN(n2627) );
  OAI22_X2 U2461 ( .A1(n419), .A2(n3186), .B1(n3185), .B2(n369), .ZN(n2628) );
  OAI22_X2 U2462 ( .A1(n419), .A2(n3187), .B1(n3186), .B2(n369), .ZN(n2629) );
  OAI22_X2 U2463 ( .A1(n419), .A2(n3188), .B1(n3187), .B2(n369), .ZN(n2630) );
  OAI22_X2 U2464 ( .A1(n419), .A2(n3189), .B1(n3188), .B2(n369), .ZN(n2631) );
  OAI22_X2 U2465 ( .A1(n419), .A2(n3190), .B1(n3189), .B2(n369), .ZN(n2632) );
  OAI22_X2 U2466 ( .A1(n419), .A2(n3191), .B1(n3190), .B2(n369), .ZN(n2633) );
  OAI22_X2 U2467 ( .A1(n419), .A2(n3192), .B1(n3191), .B2(n369), .ZN(n2634) );
  OAI22_X2 U2468 ( .A1(n419), .A2(n3193), .B1(n3192), .B2(n369), .ZN(n2635) );
  OAI22_X2 U2469 ( .A1(n419), .A2(n3194), .B1(n3193), .B2(n369), .ZN(n2636) );
  NAND2_X4 U2544 ( .A1(n3231), .A2(n3458), .ZN(n455) );
  XOR2_X2 U2545 ( .A(a[24]), .B(n357), .Z(n3231) );
  XOR2_X2 U2557 ( .A(a[16]), .B(n345), .Z(n3235) );
  NAND2_X4 U2577 ( .A1(n3242), .A2(n372), .ZN(n422) );
  XOR2_X2 U2578 ( .A(a[2]), .B(n324), .Z(n3242) );
  INV_X2 U2585 ( .A(a[20]), .ZN(n3409) );
  INV_X2 U2586 ( .A(a[20]), .ZN(n3731) );
  INV_X1 U2587 ( .A(n3455), .ZN(n3410) );
  INV_X8 U2588 ( .A(n3454), .ZN(n3455) );
  INV_X1 U2589 ( .A(n366), .ZN(n416) );
  INV_X1 U2590 ( .A(n339), .ZN(n3286) );
  INV_X1 U2591 ( .A(n339), .ZN(n3571) );
  INV_X1 U2592 ( .A(n351), .ZN(n3282) );
  INV_X1 U2593 ( .A(n351), .ZN(n3611) );
  INV_X2 U2594 ( .A(n330), .ZN(n3632) );
  XNOR2_X1 U2595 ( .A(n465), .B(n3578), .ZN(n3194) );
  XNOR2_X1 U2596 ( .A(n465), .B(n3740), .ZN(n3128) );
  AND2_X1 U2597 ( .A1(n465), .A2(n366), .ZN(n2093) );
  XNOR2_X1 U2598 ( .A(n465), .B(n3531), .ZN(n3062) );
  XNOR2_X1 U2599 ( .A(n465), .B(n3438), .ZN(n3029) );
  XNOR2_X1 U2600 ( .A(n465), .B(n324), .ZN(n3161) );
  XNOR2_X1 U2601 ( .A(n465), .B(n3712), .ZN(n2930) );
  XNOR2_X1 U2602 ( .A(n465), .B(n342), .ZN(n2963) );
  XNOR2_X1 U2603 ( .A(n465), .B(n3605), .ZN(n2831) );
  XNOR2_X1 U2604 ( .A(n465), .B(n360), .ZN(n2765) );
  XNOR2_X1 U2605 ( .A(n465), .B(n348), .ZN(n2897) );
  XNOR2_X1 U2606 ( .A(n465), .B(n330), .ZN(n3095) );
  XNOR2_X1 U2607 ( .A(n465), .B(n339), .ZN(n2996) );
  XNOR2_X1 U2608 ( .A(n465), .B(n366), .ZN(n2699) );
  XNOR2_X1 U2609 ( .A(n465), .B(n351), .ZN(n2864) );
  XNOR2_X1 U2610 ( .A(n465), .B(n363), .ZN(n2732) );
  XNOR2_X1 U2611 ( .A(n465), .B(n357), .ZN(n2798) );
  INV_X1 U2612 ( .A(n465), .ZN(n3753) );
  INV_X2 U2613 ( .A(n327), .ZN(n3478) );
  INV_X2 U2614 ( .A(a[22]), .ZN(n3610) );
  XOR2_X1 U2615 ( .A(a[26]), .B(n360), .Z(n3230) );
  INV_X2 U2616 ( .A(a[4]), .ZN(n3748) );
  INV_X2 U2617 ( .A(a[12]), .ZN(n3640) );
  INV_X4 U2618 ( .A(a[30]), .ZN(n3644) );
  INV_X2 U2619 ( .A(a[8]), .ZN(n3752) );
  INV_X2 U2620 ( .A(a[24]), .ZN(n3729) );
  INV_X1 U2621 ( .A(a[2]), .ZN(n3750) );
  NAND2_X1 U2622 ( .A1(n333), .A2(a[10]), .ZN(n3500) );
  INV_X1 U2623 ( .A(a[18]), .ZN(n3587) );
  AND2_X1 U2624 ( .A1(n465), .A2(a[0]), .ZN(product[0]) );
  OAI21_X1 U2625 ( .B1(a[0]), .B2(n3754), .A(n3578), .ZN(n2604) );
  XNOR2_X1 U2626 ( .A(n469), .B(n3578), .ZN(n3193) );
  XNOR2_X1 U2627 ( .A(n469), .B(n3531), .ZN(n3061) );
  XNOR2_X1 U2628 ( .A(n469), .B(n3740), .ZN(n3127) );
  INV_X1 U2629 ( .A(n469), .ZN(n2667) );
  XNOR2_X1 U2630 ( .A(n469), .B(n3438), .ZN(n3028) );
  XNOR2_X1 U2631 ( .A(n469), .B(n324), .ZN(n3160) );
  XNOR2_X1 U2632 ( .A(n469), .B(n330), .ZN(n3094) );
  XNOR2_X1 U2633 ( .A(n469), .B(n351), .ZN(n2863) );
  XNOR2_X1 U2634 ( .A(n469), .B(n3712), .ZN(n2929) );
  XNOR2_X1 U2635 ( .A(n469), .B(n342), .ZN(n2962) );
  XNOR2_X1 U2636 ( .A(n469), .B(n363), .ZN(n2731) );
  XNOR2_X1 U2637 ( .A(n469), .B(n366), .ZN(n2698) );
  XNOR2_X1 U2638 ( .A(n469), .B(n339), .ZN(n2995) );
  XNOR2_X1 U2639 ( .A(n469), .B(n348), .ZN(n2896) );
  XNOR2_X1 U2640 ( .A(n469), .B(n360), .ZN(n2764) );
  XNOR2_X1 U2641 ( .A(n469), .B(n357), .ZN(n2797) );
  XNOR2_X1 U2642 ( .A(n471), .B(n324), .ZN(n3159) );
  XNOR2_X1 U2643 ( .A(n471), .B(n3578), .ZN(n3192) );
  XNOR2_X1 U2644 ( .A(n471), .B(n3531), .ZN(n3060) );
  INV_X1 U2645 ( .A(n471), .ZN(n2666) );
  XNOR2_X1 U2646 ( .A(n471), .B(n3740), .ZN(n3126) );
  XNOR2_X1 U2647 ( .A(n471), .B(n3438), .ZN(n3027) );
  XNOR2_X1 U2648 ( .A(n471), .B(n330), .ZN(n3093) );
  XNOR2_X1 U2649 ( .A(n471), .B(n3712), .ZN(n2928) );
  XNOR2_X1 U2650 ( .A(n471), .B(n339), .ZN(n2994) );
  XNOR2_X1 U2651 ( .A(n471), .B(n342), .ZN(n2961) );
  XNOR2_X1 U2652 ( .A(n471), .B(n351), .ZN(n2862) );
  XNOR2_X1 U2653 ( .A(n471), .B(n366), .ZN(n2697) );
  XNOR2_X1 U2654 ( .A(n471), .B(n348), .ZN(n2895) );
  XNOR2_X1 U2655 ( .A(n471), .B(n357), .ZN(n2796) );
  XNOR2_X1 U2656 ( .A(n471), .B(n360), .ZN(n2763) );
  XNOR2_X1 U2657 ( .A(n473), .B(n324), .ZN(n3158) );
  XNOR2_X1 U2658 ( .A(n473), .B(n3531), .ZN(n3059) );
  INV_X1 U2659 ( .A(n473), .ZN(n2665) );
  XNOR2_X1 U2660 ( .A(n473), .B(n3578), .ZN(n3191) );
  XNOR2_X1 U2661 ( .A(n473), .B(n3726), .ZN(n3125) );
  XNOR2_X1 U2662 ( .A(n473), .B(n330), .ZN(n3092) );
  XNOR2_X1 U2663 ( .A(n473), .B(n363), .ZN(n2729) );
  XNOR2_X1 U2664 ( .A(n473), .B(n348), .ZN(n2894) );
  XNOR2_X1 U2665 ( .A(n473), .B(n3712), .ZN(n2927) );
  XNOR2_X1 U2666 ( .A(n473), .B(n342), .ZN(n2960) );
  XNOR2_X1 U2667 ( .A(n473), .B(n339), .ZN(n2993) );
  XNOR2_X1 U2668 ( .A(n473), .B(n357), .ZN(n2795) );
  XNOR2_X1 U2669 ( .A(n473), .B(n351), .ZN(n2861) );
  XNOR2_X1 U2670 ( .A(n473), .B(n366), .ZN(n2696) );
  XNOR2_X1 U2671 ( .A(n473), .B(n360), .ZN(n2762) );
  XNOR2_X1 U2672 ( .A(n477), .B(n330), .ZN(n3090) );
  INV_X1 U2673 ( .A(n477), .ZN(n2663) );
  XNOR2_X1 U2674 ( .A(n477), .B(n3578), .ZN(n3189) );
  XNOR2_X1 U2675 ( .A(n477), .B(n324), .ZN(n3156) );
  XNOR2_X1 U2676 ( .A(n477), .B(n3726), .ZN(n3123) );
  XNOR2_X1 U2677 ( .A(n477), .B(n339), .ZN(n2991) );
  XNOR2_X1 U2678 ( .A(n477), .B(n342), .ZN(n2958) );
  XNOR2_X1 U2679 ( .A(n477), .B(n360), .ZN(n2760) );
  XNOR2_X1 U2680 ( .A(n477), .B(n366), .ZN(n2694) );
  XNOR2_X1 U2681 ( .A(n477), .B(n363), .ZN(n2727) );
  XNOR2_X1 U2682 ( .A(n477), .B(n348), .ZN(n2892) );
  XNOR2_X1 U2683 ( .A(n477), .B(n351), .ZN(n2859) );
  XNOR2_X1 U2684 ( .A(n477), .B(n357), .ZN(n2793) );
  XNOR2_X1 U2685 ( .A(n475), .B(n3578), .ZN(n3190) );
  XNOR2_X1 U2686 ( .A(n475), .B(n324), .ZN(n3157) );
  INV_X1 U2687 ( .A(n475), .ZN(n2664) );
  XNOR2_X1 U2688 ( .A(n475), .B(n3531), .ZN(n3058) );
  XNOR2_X1 U2689 ( .A(n475), .B(n3726), .ZN(n3124) );
  XNOR2_X1 U2690 ( .A(n475), .B(n330), .ZN(n3091) );
  XNOR2_X1 U2691 ( .A(n475), .B(n339), .ZN(n2992) );
  XNOR2_X1 U2692 ( .A(n475), .B(n363), .ZN(n2728) );
  XNOR2_X1 U2693 ( .A(n475), .B(n342), .ZN(n2959) );
  XNOR2_X1 U2694 ( .A(n475), .B(n366), .ZN(n2695) );
  XNOR2_X1 U2695 ( .A(n475), .B(n3712), .ZN(n2926) );
  XNOR2_X1 U2696 ( .A(n475), .B(n348), .ZN(n2893) );
  XNOR2_X1 U2697 ( .A(n475), .B(n351), .ZN(n2860) );
  XNOR2_X1 U2698 ( .A(n475), .B(n357), .ZN(n2794) );
  XNOR2_X1 U2699 ( .A(n475), .B(n360), .ZN(n2761) );
  INV_X1 U2700 ( .A(n479), .ZN(n2662) );
  XNOR2_X1 U2701 ( .A(n479), .B(n3578), .ZN(n3188) );
  XNOR2_X1 U2702 ( .A(n479), .B(n324), .ZN(n3155) );
  XNOR2_X1 U2703 ( .A(n479), .B(n330), .ZN(n3089) );
  XNOR2_X1 U2704 ( .A(n479), .B(n3726), .ZN(n3122) );
  XNOR2_X1 U2705 ( .A(n479), .B(n339), .ZN(n2990) );
  XNOR2_X1 U2706 ( .A(n479), .B(n363), .ZN(n2726) );
  XNOR2_X1 U2707 ( .A(n479), .B(n3712), .ZN(n2924) );
  XNOR2_X1 U2708 ( .A(n479), .B(n357), .ZN(n2792) );
  XNOR2_X1 U2709 ( .A(n479), .B(n342), .ZN(n2957) );
  XNOR2_X1 U2710 ( .A(n479), .B(n348), .ZN(n2891) );
  XNOR2_X1 U2711 ( .A(n479), .B(n360), .ZN(n2759) );
  XNOR2_X1 U2712 ( .A(n479), .B(n366), .ZN(n2693) );
  XNOR2_X1 U2713 ( .A(n479), .B(n351), .ZN(n2858) );
  XNOR2_X1 U2714 ( .A(n481), .B(n3578), .ZN(n3187) );
  XNOR2_X1 U2715 ( .A(n481), .B(n330), .ZN(n3088) );
  XNOR2_X1 U2716 ( .A(n481), .B(n3438), .ZN(n3022) );
  INV_X1 U2717 ( .A(n481), .ZN(n2661) );
  XNOR2_X1 U2718 ( .A(n481), .B(n324), .ZN(n3154) );
  XNOR2_X1 U2719 ( .A(n481), .B(n3531), .ZN(n3055) );
  XNOR2_X1 U2720 ( .A(n481), .B(n357), .ZN(n2791) );
  XNOR2_X1 U2721 ( .A(n481), .B(n3726), .ZN(n3121) );
  XNOR2_X1 U2722 ( .A(n481), .B(n351), .ZN(n2857) );
  XNOR2_X1 U2723 ( .A(n481), .B(n363), .ZN(n2725) );
  XNOR2_X1 U2724 ( .A(n481), .B(n3712), .ZN(n2923) );
  XNOR2_X1 U2725 ( .A(n481), .B(n342), .ZN(n2956) );
  XNOR2_X1 U2726 ( .A(n481), .B(n339), .ZN(n2989) );
  XNOR2_X1 U2727 ( .A(n481), .B(n348), .ZN(n2890) );
  XNOR2_X1 U2728 ( .A(n481), .B(n366), .ZN(n2692) );
  INV_X1 U2729 ( .A(n485), .ZN(n2659) );
  XNOR2_X1 U2730 ( .A(n485), .B(n3726), .ZN(n3119) );
  XNOR2_X1 U2731 ( .A(n485), .B(n3578), .ZN(n3185) );
  XNOR2_X1 U2732 ( .A(n485), .B(n330), .ZN(n3086) );
  XNOR2_X1 U2733 ( .A(n485), .B(n324), .ZN(n3152) );
  XNOR2_X1 U2734 ( .A(n485), .B(n357), .ZN(n2789) );
  XNOR2_X1 U2735 ( .A(n485), .B(n360), .ZN(n2756) );
  XNOR2_X1 U2736 ( .A(n485), .B(n339), .ZN(n2987) );
  XNOR2_X1 U2737 ( .A(n485), .B(n366), .ZN(n2690) );
  XNOR2_X1 U2738 ( .A(n485), .B(n3712), .ZN(n2921) );
  XNOR2_X1 U2739 ( .A(n485), .B(n348), .ZN(n2888) );
  XNOR2_X1 U2740 ( .A(n485), .B(n351), .ZN(n2855) );
  XNOR2_X1 U2741 ( .A(n485), .B(n342), .ZN(n2954) );
  INV_X1 U2742 ( .A(n483), .ZN(n2660) );
  XNOR2_X1 U2743 ( .A(n483), .B(n3726), .ZN(n3120) );
  XNOR2_X1 U2744 ( .A(n483), .B(n3578), .ZN(n3186) );
  XNOR2_X1 U2745 ( .A(n483), .B(n330), .ZN(n3087) );
  XNOR2_X1 U2746 ( .A(n483), .B(n357), .ZN(n2790) );
  XNOR2_X1 U2747 ( .A(n483), .B(n324), .ZN(n3153) );
  XNOR2_X1 U2748 ( .A(n483), .B(n363), .ZN(n2724) );
  XNOR2_X1 U2749 ( .A(n483), .B(n342), .ZN(n2955) );
  XNOR2_X1 U2750 ( .A(n483), .B(n366), .ZN(n2691) );
  XNOR2_X1 U2751 ( .A(n483), .B(n3712), .ZN(n2922) );
  XNOR2_X1 U2752 ( .A(n483), .B(n360), .ZN(n2757) );
  XNOR2_X1 U2753 ( .A(n483), .B(n351), .ZN(n2856) );
  XNOR2_X1 U2754 ( .A(n483), .B(n348), .ZN(n2889) );
  XNOR2_X1 U2755 ( .A(n483), .B(n339), .ZN(n2988) );
  INV_X1 U2756 ( .A(n487), .ZN(n2658) );
  XNOR2_X1 U2757 ( .A(n487), .B(n324), .ZN(n3151) );
  XNOR2_X1 U2758 ( .A(n487), .B(n330), .ZN(n3085) );
  XNOR2_X1 U2759 ( .A(n487), .B(n366), .ZN(n2689) );
  XNOR2_X1 U2760 ( .A(n487), .B(n3726), .ZN(n3118) );
  XNOR2_X1 U2761 ( .A(n487), .B(n3712), .ZN(n2920) );
  XNOR2_X1 U2762 ( .A(n487), .B(n360), .ZN(n2755) );
  XNOR2_X1 U2763 ( .A(n487), .B(n357), .ZN(n2788) );
  XNOR2_X1 U2764 ( .A(n487), .B(n339), .ZN(n2986) );
  XNOR2_X1 U2765 ( .A(n487), .B(n351), .ZN(n2854) );
  XNOR2_X1 U2766 ( .A(n487), .B(n348), .ZN(n2887) );
  XNOR2_X1 U2767 ( .A(n487), .B(n342), .ZN(n2953) );
  INV_X1 U2768 ( .A(n489), .ZN(n2657) );
  XNOR2_X1 U2769 ( .A(n489), .B(n330), .ZN(n3084) );
  XNOR2_X1 U2770 ( .A(n489), .B(n366), .ZN(n2688) );
  XNOR2_X1 U2771 ( .A(n489), .B(n324), .ZN(n3150) );
  XNOR2_X1 U2772 ( .A(n489), .B(n357), .ZN(n2787) );
  XNOR2_X1 U2773 ( .A(n489), .B(n3726), .ZN(n3117) );
  XNOR2_X1 U2774 ( .A(n489), .B(n3712), .ZN(n2919) );
  XNOR2_X1 U2775 ( .A(n489), .B(n342), .ZN(n2952) );
  XNOR2_X1 U2776 ( .A(n489), .B(n360), .ZN(n2754) );
  XNOR2_X1 U2777 ( .A(n489), .B(n339), .ZN(n2985) );
  XNOR2_X1 U2778 ( .A(n489), .B(n351), .ZN(n2853) );
  XNOR2_X1 U2779 ( .A(n489), .B(n363), .ZN(n2721) );
  XNOR2_X1 U2780 ( .A(n489), .B(n348), .ZN(n2886) );
  INV_X1 U2781 ( .A(n493), .ZN(n2655) );
  XNOR2_X1 U2782 ( .A(n493), .B(n3438), .ZN(n3016) );
  XNOR2_X1 U2783 ( .A(n493), .B(n324), .ZN(n3148) );
  XNOR2_X1 U2784 ( .A(n493), .B(n351), .ZN(n2851) );
  XNOR2_X1 U2785 ( .A(n493), .B(n363), .ZN(n2719) );
  XNOR2_X1 U2786 ( .A(n493), .B(n366), .ZN(n2686) );
  XNOR2_X1 U2787 ( .A(n493), .B(n330), .ZN(n3082) );
  XNOR2_X1 U2788 ( .A(n493), .B(n357), .ZN(n2785) );
  XNOR2_X1 U2789 ( .A(n493), .B(n342), .ZN(n2950) );
  XNOR2_X1 U2790 ( .A(n493), .B(n3712), .ZN(n2917) );
  XNOR2_X1 U2791 ( .A(n493), .B(n339), .ZN(n2983) );
  XNOR2_X1 U2792 ( .A(n493), .B(n360), .ZN(n2752) );
  INV_X1 U2793 ( .A(n491), .ZN(n2656) );
  XNOR2_X1 U2794 ( .A(n491), .B(n3726), .ZN(n3116) );
  XNOR2_X1 U2795 ( .A(n491), .B(n351), .ZN(n2852) );
  XNOR2_X1 U2796 ( .A(n491), .B(n363), .ZN(n2720) );
  XNOR2_X1 U2797 ( .A(n491), .B(n357), .ZN(n2786) );
  XNOR2_X1 U2798 ( .A(n491), .B(n330), .ZN(n3083) );
  XNOR2_X1 U2799 ( .A(n491), .B(n366), .ZN(n2687) );
  XNOR2_X1 U2800 ( .A(n491), .B(n324), .ZN(n3149) );
  XNOR2_X1 U2801 ( .A(n491), .B(n342), .ZN(n2951) );
  XNOR2_X1 U2802 ( .A(n491), .B(n339), .ZN(n2984) );
  XNOR2_X1 U2803 ( .A(n491), .B(n360), .ZN(n2753) );
  XNOR2_X1 U2804 ( .A(n491), .B(n3712), .ZN(n2918) );
  INV_X1 U2805 ( .A(n495), .ZN(n2654) );
  XNOR2_X1 U2806 ( .A(n495), .B(n351), .ZN(n2850) );
  XNOR2_X1 U2807 ( .A(n495), .B(n360), .ZN(n2751) );
  XNOR2_X1 U2808 ( .A(n495), .B(n330), .ZN(n3081) );
  XNOR2_X1 U2809 ( .A(n495), .B(n363), .ZN(n2718) );
  XNOR2_X1 U2810 ( .A(n495), .B(n324), .ZN(n3147) );
  XNOR2_X1 U2811 ( .A(n495), .B(n366), .ZN(n2685) );
  XNOR2_X1 U2812 ( .A(n495), .B(n3712), .ZN(n2916) );
  XNOR2_X1 U2813 ( .A(n495), .B(n339), .ZN(n2982) );
  XNOR2_X1 U2814 ( .A(n495), .B(n357), .ZN(n2784) );
  XNOR2_X1 U2815 ( .A(n495), .B(n342), .ZN(n2949) );
  INV_X1 U2816 ( .A(n497), .ZN(n2653) );
  XNOR2_X1 U2817 ( .A(n497), .B(n324), .ZN(n3146) );
  XNOR2_X1 U2818 ( .A(n497), .B(n360), .ZN(n2750) );
  XNOR2_X1 U2819 ( .A(n497), .B(n363), .ZN(n2717) );
  XNOR2_X1 U2820 ( .A(n497), .B(n330), .ZN(n3080) );
  XNOR2_X1 U2821 ( .A(n497), .B(n357), .ZN(n2783) );
  XNOR2_X1 U2822 ( .A(n497), .B(n351), .ZN(n2849) );
  XNOR2_X1 U2823 ( .A(n497), .B(n366), .ZN(n2684) );
  XNOR2_X1 U2824 ( .A(n497), .B(n339), .ZN(n2981) );
  XNOR2_X1 U2825 ( .A(n497), .B(n3726), .ZN(n3113) );
  XNOR2_X1 U2826 ( .A(n497), .B(n342), .ZN(n2948) );
  INV_X1 U2827 ( .A(n501), .ZN(n2651) );
  XNOR2_X1 U2828 ( .A(n501), .B(n3726), .ZN(n3111) );
  XNOR2_X1 U2829 ( .A(n501), .B(n357), .ZN(n2781) );
  XNOR2_X1 U2830 ( .A(n501), .B(n330), .ZN(n3078) );
  XNOR2_X1 U2831 ( .A(n501), .B(n363), .ZN(n2715) );
  XNOR2_X1 U2832 ( .A(n501), .B(n366), .ZN(n2682) );
  XNOR2_X1 U2833 ( .A(n501), .B(n3712), .ZN(n2913) );
  XNOR2_X1 U2834 ( .A(n501), .B(n360), .ZN(n2748) );
  XNOR2_X1 U2835 ( .A(n501), .B(n351), .ZN(n2847) );
  XNOR2_X1 U2836 ( .A(n501), .B(n324), .ZN(n3144) );
  XNOR2_X1 U2837 ( .A(n501), .B(n342), .ZN(n2946) );
  XNOR2_X1 U2838 ( .A(n501), .B(n339), .ZN(n2979) );
  INV_X1 U2839 ( .A(n499), .ZN(n2652) );
  XNOR2_X1 U2840 ( .A(n499), .B(n357), .ZN(n2782) );
  XNOR2_X1 U2841 ( .A(n499), .B(n330), .ZN(n3079) );
  XNOR2_X1 U2842 ( .A(n499), .B(n360), .ZN(n2749) );
  XNOR2_X1 U2843 ( .A(n499), .B(n363), .ZN(n2716) );
  XNOR2_X1 U2844 ( .A(n499), .B(n351), .ZN(n2848) );
  XNOR2_X1 U2845 ( .A(n499), .B(n348), .ZN(n2881) );
  XNOR2_X1 U2846 ( .A(n499), .B(n3712), .ZN(n2914) );
  XNOR2_X1 U2847 ( .A(n499), .B(n324), .ZN(n3145) );
  XNOR2_X1 U2848 ( .A(n499), .B(n366), .ZN(n2683) );
  XNOR2_X1 U2849 ( .A(n499), .B(n339), .ZN(n2980) );
  XNOR2_X1 U2850 ( .A(n499), .B(n3726), .ZN(n3112) );
  XNOR2_X1 U2851 ( .A(n499), .B(n342), .ZN(n2947) );
  INV_X1 U2852 ( .A(n503), .ZN(n2650) );
  XNOR2_X1 U2853 ( .A(n503), .B(n3605), .ZN(n2813) );
  XNOR2_X1 U2854 ( .A(n503), .B(n3726), .ZN(n3110) );
  XNOR2_X1 U2855 ( .A(n503), .B(n342), .ZN(n2945) );
  XNOR2_X1 U2856 ( .A(n503), .B(n357), .ZN(n2780) );
  XNOR2_X1 U2857 ( .A(n503), .B(n366), .ZN(n2681) );
  XNOR2_X1 U2858 ( .A(n503), .B(n324), .ZN(n3143) );
  XNOR2_X1 U2859 ( .A(n503), .B(n351), .ZN(n2846) );
  XNOR2_X1 U2860 ( .A(n503), .B(n363), .ZN(n2714) );
  XNOR2_X1 U2861 ( .A(n503), .B(n3712), .ZN(n2912) );
  XNOR2_X1 U2862 ( .A(n503), .B(n360), .ZN(n2747) );
  XNOR2_X1 U2863 ( .A(n503), .B(n339), .ZN(n2978) );
  INV_X1 U2864 ( .A(n505), .ZN(n2649) );
  XNOR2_X1 U2865 ( .A(n505), .B(n3438), .ZN(n3010) );
  XNOR2_X1 U2866 ( .A(n505), .B(n366), .ZN(n2680) );
  XNOR2_X1 U2867 ( .A(n505), .B(n342), .ZN(n2944) );
  XNOR2_X1 U2868 ( .A(n505), .B(n3712), .ZN(n2911) );
  XNOR2_X1 U2869 ( .A(n505), .B(n3726), .ZN(n3109) );
  XNOR2_X1 U2870 ( .A(n505), .B(n324), .ZN(n3142) );
  XNOR2_X1 U2871 ( .A(n505), .B(n360), .ZN(n2746) );
  XNOR2_X1 U2872 ( .A(n505), .B(n357), .ZN(n2779) );
  XNOR2_X1 U2873 ( .A(n505), .B(n363), .ZN(n2713) );
  XNOR2_X1 U2874 ( .A(n505), .B(n351), .ZN(n2845) );
  XNOR2_X1 U2875 ( .A(n505), .B(n348), .ZN(n2878) );
  XNOR2_X1 U2876 ( .A(n505), .B(n339), .ZN(n2977) );
  INV_X1 U2877 ( .A(n509), .ZN(n2647) );
  XNOR2_X1 U2878 ( .A(n509), .B(n363), .ZN(n2711) );
  XNOR2_X1 U2879 ( .A(n509), .B(n330), .ZN(n3074) );
  XNOR2_X1 U2880 ( .A(n509), .B(n324), .ZN(n3140) );
  XNOR2_X1 U2881 ( .A(n509), .B(n366), .ZN(n2678) );
  XNOR2_X1 U2882 ( .A(n509), .B(n360), .ZN(n2744) );
  XNOR2_X1 U2883 ( .A(n509), .B(n3726), .ZN(n3107) );
  XNOR2_X1 U2884 ( .A(n509), .B(n351), .ZN(n2843) );
  XNOR2_X1 U2885 ( .A(n509), .B(n357), .ZN(n2777) );
  XNOR2_X1 U2886 ( .A(n509), .B(n342), .ZN(n2942) );
  XNOR2_X1 U2887 ( .A(n509), .B(n339), .ZN(n2975) );
  XNOR2_X1 U2888 ( .A(n509), .B(n348), .ZN(n2876) );
  XNOR2_X1 U2889 ( .A(n509), .B(n3712), .ZN(n2909) );
  INV_X1 U2890 ( .A(n507), .ZN(n2648) );
  XNOR2_X1 U2891 ( .A(n507), .B(n363), .ZN(n2712) );
  XNOR2_X1 U2892 ( .A(n507), .B(n366), .ZN(n2679) );
  XNOR2_X1 U2893 ( .A(n507), .B(n324), .ZN(n3141) );
  XNOR2_X1 U2894 ( .A(n507), .B(n360), .ZN(n2745) );
  XNOR2_X1 U2895 ( .A(n507), .B(n342), .ZN(n2943) );
  XNOR2_X1 U2896 ( .A(n507), .B(n339), .ZN(n2976) );
  XNOR2_X1 U2897 ( .A(n507), .B(n3726), .ZN(n3108) );
  XNOR2_X1 U2898 ( .A(n507), .B(n3712), .ZN(n2910) );
  XNOR2_X1 U2899 ( .A(n507), .B(n351), .ZN(n2844) );
  XNOR2_X1 U2900 ( .A(n507), .B(n357), .ZN(n2778) );
  XNOR2_X1 U2901 ( .A(n507), .B(n348), .ZN(n2877) );
  INV_X1 U2902 ( .A(n511), .ZN(n2646) );
  XNOR2_X1 U2903 ( .A(n511), .B(n360), .ZN(n2743) );
  XNOR2_X1 U2904 ( .A(n511), .B(n363), .ZN(n2710) );
  XNOR2_X1 U2905 ( .A(n511), .B(n348), .ZN(n2875) );
  XNOR2_X1 U2906 ( .A(n511), .B(n3438), .ZN(n3007) );
  XNOR2_X1 U2907 ( .A(n511), .B(n324), .ZN(n3139) );
  XNOR2_X1 U2908 ( .A(n511), .B(n366), .ZN(n2677) );
  XNOR2_X1 U2909 ( .A(n511), .B(n351), .ZN(n2842) );
  XNOR2_X1 U2910 ( .A(n511), .B(n357), .ZN(n2776) );
  XNOR2_X1 U2911 ( .A(n511), .B(n339), .ZN(n2974) );
  XNOR2_X1 U2912 ( .A(n511), .B(n3726), .ZN(n3106) );
  XNOR2_X1 U2913 ( .A(n511), .B(n342), .ZN(n2941) );
  XNOR2_X1 U2914 ( .A(n511), .B(n330), .ZN(n3073) );
  XNOR2_X1 U2915 ( .A(n511), .B(n3712), .ZN(n2908) );
  INV_X1 U2916 ( .A(n513), .ZN(n2645) );
  XNOR2_X1 U2917 ( .A(n513), .B(n360), .ZN(n2742) );
  XNOR2_X1 U2918 ( .A(n513), .B(n363), .ZN(n2709) );
  XNOR2_X1 U2919 ( .A(n513), .B(n342), .ZN(n2940) );
  XNOR2_X1 U2920 ( .A(n513), .B(n366), .ZN(n2676) );
  XNOR2_X1 U2921 ( .A(n513), .B(n351), .ZN(n2841) );
  XNOR2_X1 U2922 ( .A(n513), .B(n348), .ZN(n2874) );
  XNOR2_X1 U2923 ( .A(n513), .B(n357), .ZN(n2775) );
  XNOR2_X1 U2924 ( .A(n513), .B(n339), .ZN(n2973) );
  XNOR2_X1 U2925 ( .A(n513), .B(n3726), .ZN(n3105) );
  XNOR2_X1 U2926 ( .A(n513), .B(n324), .ZN(n3138) );
  XNOR2_X1 U2927 ( .A(n513), .B(n330), .ZN(n3072) );
  XNOR2_X1 U2928 ( .A(n513), .B(n3712), .ZN(n2907) );
  INV_X1 U2929 ( .A(n517), .ZN(n2643) );
  XNOR2_X1 U2930 ( .A(n517), .B(n366), .ZN(n2674) );
  XNOR2_X1 U2931 ( .A(n517), .B(n357), .ZN(n2773) );
  XNOR2_X1 U2932 ( .A(n517), .B(n363), .ZN(n2707) );
  XNOR2_X1 U2933 ( .A(n517), .B(n3712), .ZN(n2905) );
  XNOR2_X1 U2934 ( .A(n517), .B(n360), .ZN(n2740) );
  XNOR2_X1 U2935 ( .A(n517), .B(n348), .ZN(n2872) );
  XNOR2_X1 U2936 ( .A(n517), .B(n339), .ZN(n2971) );
  XNOR2_X1 U2937 ( .A(n517), .B(n330), .ZN(n3070) );
  XNOR2_X1 U2938 ( .A(n517), .B(n324), .ZN(n3136) );
  XNOR2_X1 U2939 ( .A(n517), .B(n351), .ZN(n2839) );
  XNOR2_X1 U2940 ( .A(n517), .B(n3726), .ZN(n3103) );
  XNOR2_X1 U2941 ( .A(n517), .B(n342), .ZN(n2938) );
  INV_X1 U2942 ( .A(n515), .ZN(n2644) );
  XNOR2_X1 U2943 ( .A(n515), .B(n363), .ZN(n2708) );
  XNOR2_X1 U2944 ( .A(n515), .B(n366), .ZN(n2675) );
  XNOR2_X1 U2945 ( .A(n515), .B(n3712), .ZN(n2906) );
  XNOR2_X1 U2946 ( .A(n515), .B(n357), .ZN(n2774) );
  XNOR2_X1 U2947 ( .A(n515), .B(n360), .ZN(n2741) );
  XNOR2_X1 U2948 ( .A(n515), .B(n351), .ZN(n2840) );
  XNOR2_X1 U2949 ( .A(n515), .B(n348), .ZN(n2873) );
  XNOR2_X1 U2950 ( .A(n515), .B(n330), .ZN(n3071) );
  XNOR2_X1 U2951 ( .A(n515), .B(n339), .ZN(n2972) );
  XNOR2_X1 U2952 ( .A(n515), .B(n3726), .ZN(n3104) );
  XNOR2_X1 U2953 ( .A(n515), .B(n342), .ZN(n2939) );
  XNOR2_X1 U2954 ( .A(n515), .B(n324), .ZN(n3137) );
  INV_X1 U2955 ( .A(n519), .ZN(n2642) );
  XNOR2_X1 U2956 ( .A(n519), .B(n366), .ZN(n2673) );
  XNOR2_X1 U2957 ( .A(n519), .B(n363), .ZN(n2706) );
  XNOR2_X1 U2958 ( .A(n519), .B(n357), .ZN(n2772) );
  XNOR2_X1 U2959 ( .A(n519), .B(n342), .ZN(n2937) );
  XNOR2_X1 U2960 ( .A(n519), .B(n3712), .ZN(n2904) );
  XNOR2_X1 U2961 ( .A(n519), .B(n360), .ZN(n2739) );
  XNOR2_X1 U2962 ( .A(n519), .B(n330), .ZN(n3069) );
  XNOR2_X1 U2963 ( .A(n519), .B(n348), .ZN(n2871) );
  XNOR2_X1 U2964 ( .A(n519), .B(n351), .ZN(n2838) );
  XNOR2_X1 U2965 ( .A(n519), .B(n324), .ZN(n3135) );
  XNOR2_X1 U2966 ( .A(n519), .B(n339), .ZN(n2970) );
  XNOR2_X1 U2967 ( .A(n519), .B(n3726), .ZN(n3102) );
  INV_X1 U2968 ( .A(n521), .ZN(n2641) );
  XNOR2_X1 U2969 ( .A(n521), .B(n366), .ZN(n2672) );
  XNOR2_X1 U2970 ( .A(n521), .B(n363), .ZN(n2705) );
  XNOR2_X1 U2971 ( .A(n521), .B(n357), .ZN(n2771) );
  XNOR2_X1 U2972 ( .A(n521), .B(n342), .ZN(n2936) );
  XNOR2_X1 U2973 ( .A(n521), .B(n3712), .ZN(n2903) );
  XNOR2_X1 U2974 ( .A(n521), .B(n3726), .ZN(n3101) );
  XNOR2_X1 U2975 ( .A(n521), .B(n360), .ZN(n2738) );
  XNOR2_X1 U2976 ( .A(n521), .B(n351), .ZN(n2837) );
  XNOR2_X1 U2977 ( .A(n521), .B(n348), .ZN(n2870) );
  XNOR2_X1 U2978 ( .A(n521), .B(n324), .ZN(n3134) );
  XNOR2_X1 U2979 ( .A(n521), .B(n339), .ZN(n2969) );
  INV_X1 U2980 ( .A(n523), .ZN(n2640) );
  XNOR2_X1 U2981 ( .A(n523), .B(n366), .ZN(n2671) );
  XNOR2_X1 U2982 ( .A(n523), .B(n363), .ZN(n2704) );
  XNOR2_X1 U2983 ( .A(n523), .B(n360), .ZN(n2737) );
  XNOR2_X1 U2984 ( .A(n523), .B(n3605), .ZN(n2803) );
  XNOR2_X1 U2985 ( .A(n523), .B(n339), .ZN(n2968) );
  XNOR2_X1 U2986 ( .A(n523), .B(n342), .ZN(n2935) );
  XNOR2_X1 U2987 ( .A(n523), .B(n3438), .ZN(n3001) );
  XNOR2_X1 U2988 ( .A(n523), .B(n357), .ZN(n2770) );
  XNOR2_X1 U2989 ( .A(n523), .B(n3712), .ZN(n2902) );
  XNOR2_X1 U2990 ( .A(n523), .B(n351), .ZN(n2836) );
  XNOR2_X1 U2991 ( .A(n523), .B(n348), .ZN(n2869) );
  XNOR2_X1 U2992 ( .A(n523), .B(n3482), .ZN(n3100) );
  XNOR2_X1 U2993 ( .A(n523), .B(n324), .ZN(n3133) );
  INV_X1 U2994 ( .A(n525), .ZN(n2639) );
  XNOR2_X1 U2995 ( .A(n525), .B(n366), .ZN(n2670) );
  XNOR2_X1 U2996 ( .A(n525), .B(n363), .ZN(n2703) );
  XNOR2_X1 U2997 ( .A(n525), .B(n360), .ZN(n2736) );
  XNOR2_X1 U2998 ( .A(n525), .B(n351), .ZN(n2835) );
  XNOR2_X1 U2999 ( .A(n525), .B(n3605), .ZN(n2802) );
  XNOR2_X1 U3000 ( .A(n525), .B(n3438), .ZN(n3000) );
  XNOR2_X1 U3001 ( .A(n525), .B(n339), .ZN(n2967) );
  XNOR2_X1 U3002 ( .A(n525), .B(n3712), .ZN(n2901) );
  XNOR2_X1 U3003 ( .A(n525), .B(n342), .ZN(n2934) );
  XNOR2_X1 U3004 ( .A(n525), .B(n357), .ZN(n2769) );
  XNOR2_X1 U3005 ( .A(n525), .B(n348), .ZN(n2868) );
  XNOR2_X1 U3006 ( .A(n525), .B(n330), .ZN(n3066) );
  XNOR2_X1 U3007 ( .A(n525), .B(n324), .ZN(n3132) );
  INV_X1 U3008 ( .A(n527), .ZN(n2638) );
  XNOR2_X1 U3009 ( .A(n527), .B(n366), .ZN(n2669) );
  XNOR2_X1 U3010 ( .A(n527), .B(n363), .ZN(n2702) );
  XNOR2_X1 U3011 ( .A(n527), .B(n360), .ZN(n2735) );
  XNOR2_X1 U3012 ( .A(n527), .B(n3438), .ZN(n2999) );
  XNOR2_X1 U3013 ( .A(n527), .B(n351), .ZN(n2834) );
  XNOR2_X1 U3014 ( .A(n527), .B(n357), .ZN(n2768) );
  XNOR2_X1 U3015 ( .A(n527), .B(n324), .ZN(n3131) );
  XNOR2_X1 U3016 ( .A(n527), .B(n348), .ZN(n2867) );
  XNOR2_X1 U3017 ( .A(n527), .B(n3712), .ZN(n2900) );
  XNOR2_X1 U3018 ( .A(n527), .B(n339), .ZN(n2966) );
  XNOR2_X1 U3019 ( .A(n527), .B(n342), .ZN(n2933) );
  XNOR2_X1 U3020 ( .A(n527), .B(n330), .ZN(n3065) );
  INV_X1 U3021 ( .A(n529), .ZN(n2637) );
  XNOR2_X1 U3022 ( .A(n529), .B(n366), .ZN(n2668) );
  XNOR2_X1 U3023 ( .A(n529), .B(n363), .ZN(n2701) );
  XNOR2_X1 U3024 ( .A(n529), .B(n360), .ZN(n2734) );
  XNOR2_X1 U3025 ( .A(n529), .B(n357), .ZN(n2767) );
  XNOR2_X1 U3026 ( .A(n529), .B(n348), .ZN(n2866) );
  XNOR2_X1 U3027 ( .A(n529), .B(n3605), .ZN(n2800) );
  XNOR2_X1 U3028 ( .A(n529), .B(n351), .ZN(n2833) );
  XNOR2_X1 U3029 ( .A(n529), .B(n324), .ZN(n3130) );
  XNOR2_X1 U3030 ( .A(n529), .B(n3726), .ZN(n3097) );
  XNOR2_X1 U3031 ( .A(n529), .B(n3712), .ZN(n2899) );
  XNOR2_X1 U3032 ( .A(n529), .B(n342), .ZN(n2932) );
  XNOR2_X1 U3033 ( .A(n529), .B(n339), .ZN(n2965) );
  XNOR2_X1 U3034 ( .A(n529), .B(n330), .ZN(n3064) );
  XNOR2_X1 U3035 ( .A(n477), .B(n354), .ZN(n2826) );
  XNOR2_X1 U3036 ( .A(n489), .B(n354), .ZN(n2820) );
  XNOR2_X1 U3037 ( .A(n519), .B(n354), .ZN(n2805) );
  XNOR2_X1 U3038 ( .A(n485), .B(n354), .ZN(n2822) );
  XNOR2_X1 U3039 ( .A(n487), .B(n354), .ZN(n2821) );
  XNOR2_X1 U3040 ( .A(n521), .B(n354), .ZN(n2804) );
  XNOR2_X1 U3041 ( .A(n513), .B(n354), .ZN(n2808) );
  XNOR2_X1 U3042 ( .A(n527), .B(n354), .ZN(n2801) );
  XNOR2_X1 U3043 ( .A(n483), .B(n354), .ZN(n2823) );
  XNOR2_X1 U3044 ( .A(n505), .B(n354), .ZN(n2812) );
  XNOR2_X1 U3045 ( .A(n491), .B(n354), .ZN(n2819) );
  XNOR2_X1 U3046 ( .A(n507), .B(n354), .ZN(n2811) );
  XNOR2_X1 U3047 ( .A(n469), .B(n354), .ZN(n2830) );
  XNOR2_X1 U3048 ( .A(n471), .B(n354), .ZN(n2829) );
  XNOR2_X1 U3049 ( .A(n509), .B(n354), .ZN(n2810) );
  XNOR2_X1 U3050 ( .A(n479), .B(n354), .ZN(n2825) );
  XNOR2_X1 U3051 ( .A(n515), .B(n354), .ZN(n2807) );
  XNOR2_X1 U3052 ( .A(n497), .B(n354), .ZN(n2816) );
  XNOR2_X1 U3053 ( .A(n473), .B(n354), .ZN(n2828) );
  XNOR2_X1 U3054 ( .A(n511), .B(n354), .ZN(n2809) );
  XNOR2_X1 U3055 ( .A(n481), .B(n354), .ZN(n2824) );
  XNOR2_X1 U3056 ( .A(n517), .B(n354), .ZN(n2806) );
  XNOR2_X1 U3057 ( .A(n475), .B(n354), .ZN(n2827) );
  XNOR2_X1 U3058 ( .A(n499), .B(n354), .ZN(n2815) );
  XNOR2_X1 U3059 ( .A(n501), .B(n354), .ZN(n2814) );
  XNOR2_X1 U3060 ( .A(n507), .B(n336), .ZN(n3009) );
  XNOR2_X1 U3061 ( .A(n491), .B(n336), .ZN(n3017) );
  XNOR2_X1 U3062 ( .A(n509), .B(n336), .ZN(n3008) );
  XNOR2_X1 U3063 ( .A(n479), .B(n336), .ZN(n3023) );
  XNOR2_X1 U3064 ( .A(n473), .B(n336), .ZN(n3026) );
  XNOR2_X1 U3065 ( .A(n519), .B(n336), .ZN(n3003) );
  XNOR2_X1 U3066 ( .A(n513), .B(n336), .ZN(n3006) );
  XNOR2_X1 U3067 ( .A(n477), .B(n336), .ZN(n3024) );
  XNOR2_X1 U3068 ( .A(n517), .B(n336), .ZN(n3004) );
  XNOR2_X1 U3069 ( .A(n489), .B(n336), .ZN(n3018) );
  XNOR2_X1 U3070 ( .A(n475), .B(n336), .ZN(n3025) );
  XNOR2_X1 U3071 ( .A(n495), .B(n336), .ZN(n3015) );
  XNOR2_X1 U3072 ( .A(n521), .B(n336), .ZN(n3002) );
  XNOR2_X1 U3073 ( .A(n483), .B(n336), .ZN(n3021) );
  XNOR2_X1 U3074 ( .A(n529), .B(n336), .ZN(n2998) );
  XNOR2_X1 U3075 ( .A(n515), .B(n336), .ZN(n3005) );
  XNOR2_X1 U3076 ( .A(n499), .B(n336), .ZN(n3013) );
  XNOR2_X1 U3077 ( .A(n503), .B(n336), .ZN(n3011) );
  XNOR2_X1 U3078 ( .A(n501), .B(n336), .ZN(n3012) );
  XNOR2_X1 U3079 ( .A(n497), .B(n336), .ZN(n3014) );
  XNOR2_X1 U3080 ( .A(n485), .B(n336), .ZN(n3020) );
  XNOR2_X1 U3081 ( .A(n487), .B(n336), .ZN(n3019) );
  INV_X1 U3082 ( .A(n336), .ZN(n3437) );
  NAND2_X1 U3083 ( .A1(n3640), .A2(n336), .ZN(n3643) );
  XOR2_X1 U3084 ( .A(a[10]), .B(n336), .Z(n3238) );
  INV_X1 U3085 ( .A(n336), .ZN(n3641) );
  BUF_X8 U3086 ( .A(n333), .Z(n3411) );
  XOR2_X1 U3087 ( .A(n1676), .B(n1678), .Z(n3412) );
  XOR2_X1 U3088 ( .A(n1701), .B(n3412), .Z(n1672) );
  NAND2_X1 U3089 ( .A1(n1701), .A2(n1676), .ZN(n3413) );
  NAND2_X1 U3090 ( .A1(n1701), .A2(n1678), .ZN(n3414) );
  NAND2_X1 U3091 ( .A1(n1676), .A2(n1678), .ZN(n3415) );
  NAND3_X1 U3092 ( .A1(n3413), .A2(n3415), .A3(n3414), .ZN(n1671) );
  OAI22_X1 U3093 ( .A1(n449), .A2(n2839), .B1(n2838), .B2(n399), .ZN(n2271) );
  AOI21_X1 U3094 ( .B1(n694), .B2(n703), .A(n695), .ZN(n693) );
  NOR2_X2 U3095 ( .A1(n699), .A2(n696), .ZN(n694) );
  NAND2_X2 U3096 ( .A1(n694), .A2(n994), .ZN(n692) );
  XOR2_X2 U3097 ( .A(n3426), .B(n1306), .Z(n1283) );
  INV_X1 U3098 ( .A(n752), .ZN(n750) );
  BUF_X1 U3099 ( .A(n1304), .Z(n3416) );
  XNOR2_X1 U3100 ( .A(n1554), .B(n3417), .ZN(n1521) );
  XNOR2_X1 U3101 ( .A(n1525), .B(n1556), .ZN(n3417) );
  XNOR2_X1 U3102 ( .A(n1495), .B(n3418), .ZN(n1491) );
  XNOR2_X1 U3103 ( .A(n1522), .B(n1524), .ZN(n3418) );
  OAI22_X1 U3104 ( .A1(n464), .A2(n2699), .B1(n2698), .B2(n3526), .ZN(n2126)
         );
  XOR2_X1 U3105 ( .A(n2407), .B(n2375), .Z(n3419) );
  XOR2_X1 U3106 ( .A(n2151), .B(n3419), .Z(n1423) );
  NAND2_X1 U3107 ( .A1(n2151), .A2(n2407), .ZN(n3420) );
  NAND2_X1 U3108 ( .A1(n2151), .A2(n2375), .ZN(n3421) );
  NAND2_X1 U3109 ( .A1(n2407), .A2(n2375), .ZN(n3422) );
  NAND3_X1 U3110 ( .A1(n3420), .A2(n3422), .A3(n3421), .ZN(n1422) );
  OR2_X1 U3111 ( .A1(n3476), .A2(n2723), .ZN(n3423) );
  OR2_X1 U3112 ( .A1(n2722), .A2(n3607), .ZN(n3424) );
  NAND2_X1 U3113 ( .A1(n3423), .A2(n3424), .ZN(n2151) );
  OAI22_X1 U3114 ( .A1(n3435), .A2(n2971), .B1(n2970), .B2(n387), .ZN(n2407)
         );
  OAI22_X1 U3115 ( .A1(n440), .A2(n2940), .B1(n2939), .B2(n390), .ZN(n2375) );
  XNOR2_X1 U3116 ( .A(n485), .B(n363), .ZN(n2723) );
  XNOR2_X1 U3117 ( .A(n487), .B(n363), .ZN(n2722) );
  INV_X1 U3118 ( .A(n753), .ZN(n751) );
  NAND2_X2 U3119 ( .A1(n3235), .A2(n3555), .ZN(n443) );
  INV_X4 U3120 ( .A(n3749), .ZN(n3425) );
  INV_X1 U3121 ( .A(n3749), .ZN(n372) );
  XNOR2_X1 U3122 ( .A(n529), .B(n321), .ZN(n3163) );
  XNOR2_X1 U3123 ( .A(n527), .B(n321), .ZN(n3164) );
  XNOR2_X1 U3124 ( .A(n525), .B(n321), .ZN(n3165) );
  XNOR2_X1 U3125 ( .A(n523), .B(n321), .ZN(n3166) );
  XNOR2_X1 U3126 ( .A(n521), .B(n321), .ZN(n3167) );
  XNOR2_X1 U3127 ( .A(n519), .B(n321), .ZN(n3168) );
  XNOR2_X1 U3128 ( .A(n517), .B(n321), .ZN(n3169) );
  XNOR2_X1 U3129 ( .A(n515), .B(n321), .ZN(n3170) );
  XNOR2_X1 U3130 ( .A(n513), .B(n321), .ZN(n3171) );
  XNOR2_X1 U3131 ( .A(n511), .B(n321), .ZN(n3172) );
  XNOR2_X1 U3132 ( .A(n509), .B(n321), .ZN(n3173) );
  XNOR2_X1 U3133 ( .A(n487), .B(n321), .ZN(n3184) );
  XNOR2_X1 U3134 ( .A(n489), .B(n321), .ZN(n3183) );
  XNOR2_X1 U3135 ( .A(n491), .B(n321), .ZN(n3182) );
  XNOR2_X1 U3136 ( .A(n493), .B(n321), .ZN(n3181) );
  XNOR2_X1 U3137 ( .A(n495), .B(n321), .ZN(n3180) );
  XNOR2_X1 U3138 ( .A(n497), .B(n321), .ZN(n3179) );
  XNOR2_X1 U3139 ( .A(n499), .B(n321), .ZN(n3178) );
  XNOR2_X1 U3140 ( .A(n501), .B(n321), .ZN(n3177) );
  XNOR2_X1 U3141 ( .A(n503), .B(n321), .ZN(n3176) );
  XNOR2_X1 U3142 ( .A(n505), .B(n321), .ZN(n3175) );
  XNOR2_X1 U3143 ( .A(n507), .B(n321), .ZN(n3174) );
  INV_X2 U3144 ( .A(n321), .ZN(n3577) );
  XNOR2_X1 U3145 ( .A(n3610), .B(n354), .ZN(n3232) );
  AOI21_X1 U3146 ( .B1(n914), .B2(n905), .A(n906), .ZN(n904) );
  OAI21_X1 U3147 ( .B1(n877), .B2(n857), .A(n858), .ZN(n856) );
  AOI21_X2 U3148 ( .B1(n906), .B2(n900), .A(n901), .ZN(n899) );
  AND2_X2 U3149 ( .A1(n3234), .A2(n3513), .ZN(n3690) );
  XOR2_X1 U3150 ( .A(n1287), .B(n1308), .Z(n3426) );
  XOR2_X1 U3151 ( .A(n1304), .B(n1285), .Z(n3427) );
  XOR2_X1 U3152 ( .A(n3427), .B(n1283), .Z(n1281) );
  NAND2_X1 U3153 ( .A1(n1287), .A2(n1308), .ZN(n3428) );
  NAND2_X1 U3154 ( .A1(n1287), .A2(n1306), .ZN(n3429) );
  NAND2_X1 U3155 ( .A1(n1308), .A2(n1306), .ZN(n3430) );
  NAND3_X1 U3156 ( .A1(n3428), .A2(n3429), .A3(n3430), .ZN(n1282) );
  NAND2_X1 U3157 ( .A1(n3416), .A2(n1285), .ZN(n3431) );
  NAND2_X1 U3158 ( .A1(n1304), .A2(n1283), .ZN(n3432) );
  NAND2_X1 U3159 ( .A1(n1285), .A2(n1283), .ZN(n3433) );
  NAND3_X1 U3160 ( .A1(n3431), .A2(n3432), .A3(n3433), .ZN(n1280) );
  INV_X1 U3161 ( .A(n3530), .ZN(n3531) );
  AOI21_X2 U3162 ( .B1(n844), .B2(n852), .A(n845), .ZN(n3434) );
  AOI21_X1 U3163 ( .B1(n844), .B2(n852), .A(n845), .ZN(n843) );
  INV_X2 U3164 ( .A(n730), .ZN(n3442) );
  XNOR2_X1 U3165 ( .A(n3570), .B(n3285), .ZN(n3236) );
  INV_X4 U3166 ( .A(n342), .ZN(n3285) );
  NAND2_X1 U3167 ( .A1(n1698), .A2(n1723), .ZN(n825) );
  NOR2_X1 U3168 ( .A1(n1698), .A2(n1723), .ZN(n824) );
  OAI22_X1 U3169 ( .A1(n464), .A2(n2691), .B1(n2690), .B2(n3526), .ZN(n2118)
         );
  AND2_X2 U3170 ( .A1(n3232), .A2(n3561), .ZN(n3676) );
  INV_X2 U3171 ( .A(n3457), .ZN(n3459) );
  OAI22_X1 U3172 ( .A1(n449), .A2(n2860), .B1(n2859), .B2(n399), .ZN(n2292) );
  INV_X4 U3173 ( .A(n3724), .ZN(n3436) );
  INV_X4 U3174 ( .A(n3724), .ZN(n3435) );
  INV_X2 U3175 ( .A(n3437), .ZN(n3438) );
  INV_X1 U3176 ( .A(n3724), .ZN(n437) );
  INV_X2 U3177 ( .A(n3753), .ZN(n3439) );
  INV_X8 U3178 ( .A(n3439), .ZN(n3440) );
  INV_X1 U3179 ( .A(n3691), .ZN(n378) );
  XOR2_X1 U3180 ( .A(n2188), .B(n2124), .Z(n3514) );
  NAND2_X1 U3181 ( .A1(n2124), .A2(n2348), .ZN(n3518) );
  OAI22_X1 U3182 ( .A1(n3477), .A2(n2702), .B1(n2701), .B2(n3557), .ZN(n2130)
         );
  OAI22_X1 U3183 ( .A1(n3477), .A2(n2705), .B1(n2704), .B2(n3557), .ZN(n2133)
         );
  OAI22_X1 U3184 ( .A1(n3477), .A2(n2709), .B1(n2708), .B2(n3557), .ZN(n2137)
         );
  OAI22_X1 U3185 ( .A1(n3477), .A2(n2708), .B1(n2707), .B2(n3557), .ZN(n2136)
         );
  OAI22_X1 U3186 ( .A1(n3477), .A2(n2711), .B1(n2710), .B2(n3557), .ZN(n2139)
         );
  OAI22_X1 U3187 ( .A1(n3477), .A2(n2707), .B1(n2706), .B2(n3557), .ZN(n2135)
         );
  OAI22_X1 U3188 ( .A1(n3477), .A2(n2713), .B1(n2712), .B2(n3557), .ZN(n2141)
         );
  OAI22_X1 U3189 ( .A1(n3477), .A2(n2710), .B1(n2709), .B2(n3557), .ZN(n2138)
         );
  OAI22_X1 U3190 ( .A1(n3477), .A2(n2725), .B1(n2724), .B2(n3557), .ZN(n2153)
         );
  OAI22_X1 U3191 ( .A1(n3477), .A2(n2715), .B1(n2714), .B2(n3557), .ZN(n2143)
         );
  OAI22_X1 U3192 ( .A1(n3477), .A2(n2720), .B1(n2719), .B2(n3557), .ZN(n2148)
         );
  OAI22_X1 U3193 ( .A1(n3477), .A2(n2730), .B1(n2729), .B2(n3557), .ZN(n2158)
         );
  NAND2_X1 U3194 ( .A1(n753), .A2(n3474), .ZN(n3441) );
  AND2_X2 U3195 ( .A1(n3441), .A2(n3442), .ZN(n3654) );
  OAI21_X2 U3196 ( .B1(n3445), .B2(n760), .A(n755), .ZN(n753) );
  NAND2_X1 U3197 ( .A1(n1011), .A2(n815), .ZN(n565) );
  AOI21_X1 U3198 ( .B1(n3497), .B2(n828), .A(n829), .ZN(n3443) );
  AOI21_X1 U3199 ( .B1(n856), .B2(n828), .A(n829), .ZN(n827) );
  NAND2_X1 U3200 ( .A1(n1012), .A2(n820), .ZN(n566) );
  XNOR2_X1 U3201 ( .A(n3644), .B(n366), .ZN(n3228) );
  OAI21_X1 U3202 ( .B1(n3670), .B2(n684), .A(n685), .ZN(n683) );
  XNOR2_X1 U3203 ( .A(n3409), .B(n351), .ZN(n3233) );
  NAND2_X1 U3204 ( .A1(n1642), .A2(n1669), .ZN(n815) );
  NAND2_X2 U3205 ( .A1(n1882), .A2(n1899), .ZN(n875) );
  NOR2_X1 U3206 ( .A1(n1882), .A2(n1899), .ZN(n874) );
  XOR2_X1 U3207 ( .A(n1644), .B(n3547), .Z(n1642) );
  OR2_X2 U3208 ( .A1(n3713), .A2(n3714), .ZN(n2249) );
  INV_X8 U3209 ( .A(n3676), .ZN(n3671) );
  INV_X2 U3210 ( .A(n3728), .ZN(n405) );
  INV_X1 U3211 ( .A(n3605), .ZN(n3281) );
  OAI22_X1 U3212 ( .A1(n3671), .A2(n2812), .B1(n2811), .B2(n402), .ZN(n2243)
         );
  XNOR2_X1 U3213 ( .A(n3640), .B(n339), .ZN(n3237) );
  OAI21_X1 U3214 ( .B1(n861), .B2(n865), .A(n862), .ZN(n860) );
  OAI21_X1 U3215 ( .B1(n3434), .B2(n830), .A(n831), .ZN(n3444) );
  OAI21_X1 U3216 ( .B1(n843), .B2(n830), .A(n831), .ZN(n829) );
  OAI21_X1 U3217 ( .B1(n855), .B2(n849), .A(n850), .ZN(n848) );
  NAND2_X1 U3218 ( .A1(n851), .A2(n850), .ZN(n571) );
  NOR2_X2 U3219 ( .A1(n1327), .A2(n1350), .ZN(n3445) );
  NOR2_X1 U3220 ( .A1(n1327), .A2(n1350), .ZN(n754) );
  OAI21_X1 U3221 ( .B1(n819), .B2(n825), .A(n820), .ZN(n3446) );
  OAI21_X1 U3222 ( .B1(n819), .B2(n825), .A(n820), .ZN(n818) );
  INV_X1 U3223 ( .A(n850), .ZN(n852) );
  OAI22_X1 U3224 ( .A1(n419), .A2(n3165), .B1(n3164), .B2(n369), .ZN(n3447) );
  OAI21_X2 U3225 ( .B1(n701), .B2(n699), .A(n700), .ZN(n698) );
  NAND2_X2 U3226 ( .A1(n832), .A2(n3480), .ZN(n830) );
  OAI22_X1 U3227 ( .A1(n437), .A2(n2984), .B1(n2983), .B2(n387), .ZN(n2420) );
  INV_X8 U3228 ( .A(n3568), .ZN(n384) );
  INV_X2 U3229 ( .A(n3533), .ZN(n3568) );
  OAI21_X1 U3230 ( .B1(n3670), .B2(n707), .A(n708), .ZN(n706) );
  NOR2_X4 U3231 ( .A1(n3449), .A2(n3747), .ZN(n3448) );
  XNOR2_X1 U3232 ( .A(a[4]), .B(n3479), .ZN(n3449) );
  NAND2_X1 U3233 ( .A1(n1554), .A2(n1525), .ZN(n3450) );
  NAND2_X2 U3234 ( .A1(n1554), .A2(n1556), .ZN(n3451) );
  NAND2_X1 U3235 ( .A1(n1525), .A2(n1556), .ZN(n3452) );
  NAND3_X1 U3236 ( .A1(n3450), .A2(n3452), .A3(n3451), .ZN(n1520) );
  INV_X1 U3237 ( .A(n3687), .ZN(n3453) );
  NAND2_X1 U3238 ( .A1(n3598), .A2(n3599), .ZN(n3687) );
  INV_X2 U3239 ( .A(n416), .ZN(n3454) );
  AOI21_X2 U3240 ( .B1(n726), .B2(n709), .A(n710), .ZN(n708) );
  AND2_X2 U3241 ( .A1(n3236), .A2(n3536), .ZN(n3622) );
  NOR2_X2 U3242 ( .A1(n861), .A2(n864), .ZN(n859) );
  NOR2_X2 U3243 ( .A1(n1820), .A2(n1841), .ZN(n861) );
  OAI21_X1 U3244 ( .B1(n785), .B2(n765), .A(n766), .ZN(n3534) );
  INV_X1 U3245 ( .A(n838), .ZN(n3456) );
  NAND2_X2 U3246 ( .A1(n1123), .A2(n1136), .ZN(n669) );
  NOR2_X1 U3247 ( .A1(n1123), .A2(n1136), .ZN(n668) );
  AOI21_X2 U3248 ( .B1(n635), .B2(n676), .A(n636), .ZN(n634) );
  OAI21_X1 U3249 ( .B1(n634), .B2(n617), .A(n618), .ZN(n616) );
  INV_X1 U3250 ( .A(n634), .ZN(n632) );
  NAND2_X2 U3251 ( .A1(n3231), .A2(n3458), .ZN(n3603) );
  NAND2_X2 U3252 ( .A1(n3231), .A2(n3458), .ZN(n3602) );
  INV_X2 U3253 ( .A(n405), .ZN(n3457) );
  INV_X1 U3254 ( .A(n3457), .ZN(n3458) );
  INV_X2 U3255 ( .A(n3457), .ZN(n3460) );
  BUF_X1 U3256 ( .A(n798), .Z(n3461) );
  XNOR2_X1 U3257 ( .A(n623), .B(n536), .ZN(product[59]) );
  NAND2_X2 U3258 ( .A1(n1842), .A2(n1861), .ZN(n865) );
  NOR2_X2 U3259 ( .A1(n3463), .A2(n3751), .ZN(n3462) );
  XNOR2_X1 U3260 ( .A(a[8]), .B(n333), .ZN(n3463) );
  NAND2_X4 U3261 ( .A1(n3633), .A2(n3634), .ZN(n3751) );
  XOR2_X1 U3262 ( .A(n1935), .B(n1922), .Z(n3464) );
  XOR2_X1 U3263 ( .A(n1920), .B(n3464), .Z(n1918) );
  NAND2_X1 U3264 ( .A1(n1920), .A2(n1935), .ZN(n3465) );
  NAND2_X1 U3265 ( .A1(n1920), .A2(n1922), .ZN(n3466) );
  NAND2_X1 U3266 ( .A1(n1935), .A2(n1922), .ZN(n3467) );
  NAND3_X1 U3267 ( .A1(n3465), .A2(n3467), .A3(n3466), .ZN(n1917) );
  BUF_X1 U3268 ( .A(n877), .Z(n3468) );
  OR2_X1 U3269 ( .A1(n3539), .A2(n3115), .ZN(n3469) );
  OR2_X1 U3270 ( .A1(n3114), .A2(n375), .ZN(n3470) );
  NAND2_X1 U3271 ( .A1(n3469), .A2(n3470), .ZN(n2555) );
  NAND2_X1 U3272 ( .A1(n1900), .A2(n1917), .ZN(n881) );
  NOR2_X1 U3273 ( .A1(n1918), .A2(n1933), .ZN(n887) );
  XNOR2_X1 U3274 ( .A(n493), .B(n3726), .ZN(n3115) );
  XNOR2_X1 U3275 ( .A(n495), .B(n3726), .ZN(n3114) );
  INV_X1 U3276 ( .A(n847), .ZN(n845) );
  OAI22_X1 U3277 ( .A1(n3576), .A2(n3615), .B1(n3162), .B2(n3425), .ZN(n2075)
         );
  OAI22_X1 U3278 ( .A1(n3576), .A2(n3160), .B1(n3159), .B2(n3425), .ZN(n2601)
         );
  OAI22_X1 U3279 ( .A1(n3576), .A2(n3157), .B1(n3156), .B2(n3425), .ZN(n2598)
         );
  OAI22_X1 U3280 ( .A1(n422), .A2(n3153), .B1(n3152), .B2(n3425), .ZN(n2594)
         );
  OAI22_X1 U3281 ( .A1(n422), .A2(n3152), .B1(n3151), .B2(n3425), .ZN(n2593)
         );
  OAI22_X1 U3282 ( .A1(n422), .A2(n3150), .B1(n3149), .B2(n3425), .ZN(n2591)
         );
  OAI22_X1 U3283 ( .A1(n3576), .A2(n3149), .B1(n3148), .B2(n3425), .ZN(n2590)
         );
  OAI22_X1 U3284 ( .A1(n422), .A2(n3140), .B1(n3139), .B2(n3425), .ZN(n2581)
         );
  OAI22_X1 U3285 ( .A1(n3576), .A2(n3146), .B1(n3145), .B2(n3425), .ZN(n2587)
         );
  OAI22_X1 U3286 ( .A1(n3575), .A2(n3138), .B1(n3137), .B2(n372), .ZN(n2579)
         );
  XNOR2_X1 U3287 ( .A(n1405), .B(n3471), .ZN(n1403) );
  XNOR2_X1 U3288 ( .A(n1432), .B(n1407), .ZN(n3471) );
  NOR2_X1 U3289 ( .A1(n1377), .A2(n1402), .ZN(n769) );
  NOR2_X1 U3290 ( .A1(n1403), .A2(n1430), .ZN(n772) );
  NAND2_X2 U3291 ( .A1(n3635), .A2(n357), .ZN(n3598) );
  AOI21_X2 U3292 ( .B1(n612), .B2(n981), .A(n607), .ZN(n605) );
  INV_X1 U3293 ( .A(n3556), .ZN(n3745) );
  INV_X1 U3294 ( .A(n3462), .ZN(n3659) );
  INV_X1 U3295 ( .A(n3478), .ZN(n3472) );
  INV_X1 U3296 ( .A(n378), .ZN(n3636) );
  NAND2_X1 U3297 ( .A1(n1862), .A2(n1881), .ZN(n870) );
  AND2_X2 U3298 ( .A1(n3735), .A2(n3736), .ZN(n831) );
  BUF_X1 U3299 ( .A(n819), .Z(n3473) );
  BUF_X4 U3300 ( .A(a[6]), .Z(n3718) );
  NOR2_X1 U3301 ( .A1(n731), .A2(n747), .ZN(n3475) );
  NOR2_X1 U3302 ( .A1(n731), .A2(n747), .ZN(n3474) );
  INV_X4 U3303 ( .A(n3674), .ZN(n3477) );
  INV_X4 U3304 ( .A(n3674), .ZN(n3476) );
  NOR2_X1 U3305 ( .A1(n731), .A2(n747), .ZN(n729) );
  INV_X1 U3306 ( .A(n3674), .ZN(n461) );
  AND2_X4 U3307 ( .A1(n3229), .A2(n3607), .ZN(n3674) );
  OAI22_X1 U3308 ( .A1(n458), .A2(n3279), .B1(n2766), .B2(n408), .ZN(n2063) );
  OAI22_X1 U3309 ( .A1(n458), .A2(n2745), .B1(n2744), .B2(n408), .ZN(n2174) );
  OAI22_X1 U3310 ( .A1(n458), .A2(n2760), .B1(n2759), .B2(n408), .ZN(n2189) );
  OAI22_X1 U3311 ( .A1(n458), .A2(n2739), .B1(n2738), .B2(n408), .ZN(n2168) );
  OAI22_X1 U3312 ( .A1(n458), .A2(n2756), .B1(n2755), .B2(n408), .ZN(n2185) );
  OAI22_X1 U3313 ( .A1(n458), .A2(n2758), .B1(n2757), .B2(n408), .ZN(n2187) );
  OAI22_X1 U3314 ( .A1(n458), .A2(n2755), .B1(n2754), .B2(n408), .ZN(n2184) );
  OAI22_X1 U3315 ( .A1(n458), .A2(n2746), .B1(n2745), .B2(n408), .ZN(n2175) );
  OR2_X1 U3316 ( .A1(n458), .A2(n2759), .ZN(n3522) );
  OAI22_X1 U3317 ( .A1(n458), .A2(n2761), .B1(n2760), .B2(n408), .ZN(n2190) );
  OAI22_X1 U3318 ( .A1(n458), .A2(n2764), .B1(n2763), .B2(n408), .ZN(n2193) );
  OAI22_X1 U3319 ( .A1(n458), .A2(n2748), .B1(n2747), .B2(n408), .ZN(n2177) );
  OAI22_X1 U3320 ( .A1(n458), .A2(n2762), .B1(n2761), .B2(n408), .ZN(n2191) );
  OAI22_X1 U3321 ( .A1(n458), .A2(n2754), .B1(n2753), .B2(n408), .ZN(n2183) );
  OAI22_X1 U3322 ( .A1(n458), .A2(n2753), .B1(n2752), .B2(n408), .ZN(n2182) );
  INV_X1 U3323 ( .A(n3478), .ZN(n3479) );
  OAI22_X1 U3324 ( .A1(n3538), .A2(n3116), .B1(n3115), .B2(n375), .ZN(n2556)
         );
  OAI22_X1 U3325 ( .A1(n3538), .A2(n3290), .B1(n3129), .B2(n375), .ZN(n2074)
         );
  OAI22_X1 U3326 ( .A1(n3538), .A2(n3125), .B1(n3124), .B2(n375), .ZN(n2565)
         );
  OAI22_X1 U3327 ( .A1(n3538), .A2(n3124), .B1(n3123), .B2(n375), .ZN(n2564)
         );
  OAI22_X1 U3328 ( .A1(n3538), .A2(n3119), .B1(n3118), .B2(n375), .ZN(n2559)
         );
  OAI22_X1 U3329 ( .A1(n3538), .A2(n3105), .B1(n3104), .B2(n375), .ZN(n2545)
         );
  OAI22_X1 U3330 ( .A1(n3538), .A2(n3120), .B1(n3119), .B2(n375), .ZN(n2560)
         );
  OAI22_X1 U3331 ( .A1(n3538), .A2(n3122), .B1(n3121), .B2(n375), .ZN(n2562)
         );
  OAI22_X1 U3332 ( .A1(n3538), .A2(n3108), .B1(n3107), .B2(n375), .ZN(n2548)
         );
  OAI22_X1 U3333 ( .A1(n3538), .A2(n3101), .B1(n3100), .B2(n375), .ZN(n2541)
         );
  OAI22_X1 U3334 ( .A1(n3538), .A2(n3106), .B1(n3105), .B2(n375), .ZN(n2546)
         );
  OAI22_X1 U3335 ( .A1(n3538), .A2(n3107), .B1(n3106), .B2(n375), .ZN(n2547)
         );
  OAI22_X1 U3336 ( .A1(n3538), .A2(n3111), .B1(n3110), .B2(n375), .ZN(n2551)
         );
  OAI22_X1 U3337 ( .A1(n3538), .A2(n3110), .B1(n3109), .B2(n375), .ZN(n2550)
         );
  OAI22_X1 U3338 ( .A1(n3538), .A2(n3098), .B1(n3097), .B2(n375), .ZN(n2538)
         );
  OR2_X2 U3339 ( .A1(n1750), .A2(n1773), .ZN(n3480) );
  INV_X1 U3340 ( .A(n3473), .ZN(n1012) );
  OAI22_X1 U3341 ( .A1(n3603), .A2(n2768), .B1(n2767), .B2(n3459), .ZN(n2198)
         );
  OAI22_X1 U3342 ( .A1(n3603), .A2(n2773), .B1(n2772), .B2(n3459), .ZN(n2203)
         );
  OAI22_X1 U3343 ( .A1(n3602), .A2(n2781), .B1(n2780), .B2(n3459), .ZN(n2211)
         );
  OAI22_X1 U3344 ( .A1(n3603), .A2(n2786), .B1(n2785), .B2(n3460), .ZN(n2216)
         );
  OAI22_X1 U3345 ( .A1(n3603), .A2(n2772), .B1(n2771), .B2(n3459), .ZN(n2202)
         );
  OAI22_X1 U3346 ( .A1(n3602), .A2(n2793), .B1(n2792), .B2(n3460), .ZN(n2223)
         );
  OAI22_X1 U3347 ( .A1(n3603), .A2(n2789), .B1(n2788), .B2(n3459), .ZN(n2219)
         );
  OAI22_X1 U3348 ( .A1(n455), .A2(n2796), .B1(n2795), .B2(n3460), .ZN(n2226)
         );
  OAI22_X1 U3349 ( .A1(n3602), .A2(n2770), .B1(n2769), .B2(n3460), .ZN(n2200)
         );
  OAI22_X1 U3350 ( .A1(n455), .A2(n2785), .B1(n2784), .B2(n3460), .ZN(n2215)
         );
  NOR2_X1 U3351 ( .A1(n1351), .A2(n1376), .ZN(n759) );
  BUF_X1 U3352 ( .A(n3495), .Z(n3481) );
  INV_X1 U3353 ( .A(n3739), .ZN(n3482) );
  INV_X1 U3354 ( .A(n3726), .ZN(n3739) );
  OAI22_X1 U3355 ( .A1(n455), .A2(n2794), .B1(n2793), .B2(n3460), .ZN(n2224)
         );
  NAND2_X1 U3356 ( .A1(n1006), .A2(n789), .ZN(n560) );
  NAND2_X1 U3357 ( .A1(n859), .A2(n868), .ZN(n3483) );
  INV_X1 U3358 ( .A(n860), .ZN(n3484) );
  AND2_X2 U3359 ( .A1(n3483), .A2(n3484), .ZN(n858) );
  XNOR2_X1 U3360 ( .A(n717), .B(n549), .ZN(product[46]) );
  NOR2_X1 U3361 ( .A1(n3638), .A2(n3440), .ZN(n2535) );
  OAI22_X1 U3362 ( .A1(n3541), .A2(n3093), .B1(n3092), .B2(n3638), .ZN(n2532)
         );
  OAI22_X1 U3363 ( .A1(n3541), .A2(n3090), .B1(n3089), .B2(n3638), .ZN(n2529)
         );
  OAI22_X1 U3364 ( .A1(n3541), .A2(n3092), .B1(n3091), .B2(n3638), .ZN(n2531)
         );
  OAI22_X1 U3365 ( .A1(n3541), .A2(n3085), .B1(n3084), .B2(n3638), .ZN(n2524)
         );
  OAI22_X1 U3366 ( .A1(n3541), .A2(n3082), .B1(n3081), .B2(n3638), .ZN(n2521)
         );
  OAI22_X1 U3367 ( .A1(n3541), .A2(n3089), .B1(n3088), .B2(n3638), .ZN(n2528)
         );
  OAI22_X1 U3368 ( .A1(n3541), .A2(n3072), .B1(n3071), .B2(n3638), .ZN(n2511)
         );
  OAI22_X1 U3369 ( .A1(n3541), .A2(n3070), .B1(n3069), .B2(n3638), .ZN(n2509)
         );
  OAI22_X1 U3370 ( .A1(n3541), .A2(n3080), .B1(n3079), .B2(n3638), .ZN(n2519)
         );
  OAI22_X1 U3371 ( .A1(n428), .A2(n3066), .B1(n3065), .B2(n3639), .ZN(n2505)
         );
  OAI22_X1 U3372 ( .A1(n428), .A2(n3064), .B1(n3639), .B2(n3632), .ZN(n2503)
         );
  NOR2_X2 U3373 ( .A1(n1670), .A2(n1697), .ZN(n819) );
  AND2_X1 U3374 ( .A1(n752), .A2(n3474), .ZN(n3485) );
  NAND2_X1 U3375 ( .A1(n360), .A2(n3656), .ZN(n3488) );
  NAND2_X1 U3376 ( .A1(n3486), .A2(n3487), .ZN(n3489) );
  NAND2_X1 U3377 ( .A1(n3488), .A2(n3489), .ZN(n3725) );
  INV_X1 U3378 ( .A(n360), .ZN(n3486) );
  INV_X1 U3379 ( .A(n3656), .ZN(n3487) );
  NOR2_X2 U3380 ( .A1(n759), .A2(n754), .ZN(n752) );
  XOR2_X1 U3381 ( .A(a[28]), .B(n363), .Z(n3229) );
  BUF_X1 U3382 ( .A(n3699), .Z(n3490) );
  NAND2_X2 U3383 ( .A1(n3748), .A2(n324), .ZN(n3616) );
  NAND2_X1 U3384 ( .A1(n752), .A2(n729), .ZN(n727) );
  NAND2_X1 U3385 ( .A1(n1495), .A2(n1522), .ZN(n3491) );
  NAND2_X1 U3386 ( .A1(n1495), .A2(n1524), .ZN(n3492) );
  NAND2_X1 U3387 ( .A1(n1522), .A2(n1524), .ZN(n3493) );
  NAND3_X1 U3388 ( .A1(n3491), .A2(n3493), .A3(n3492), .ZN(n1490) );
  NAND2_X2 U3389 ( .A1(n3242), .A2(n372), .ZN(n3575) );
  OAI22_X1 U3390 ( .A1(n3575), .A2(n3134), .B1(n3133), .B2(n3425), .ZN(n2575)
         );
  OAI22_X1 U3391 ( .A1(n3576), .A2(n3131), .B1(n3130), .B2(n3425), .ZN(n2572)
         );
  OAI22_X1 U3392 ( .A1(n422), .A2(n3142), .B1(n3141), .B2(n3425), .ZN(n2583)
         );
  OAI22_X1 U3393 ( .A1(n3576), .A2(n3151), .B1(n3150), .B2(n3425), .ZN(n2592)
         );
  OAI22_X1 U3394 ( .A1(n3576), .A2(n3158), .B1(n3157), .B2(n3425), .ZN(n2599)
         );
  OAI22_X1 U3395 ( .A1(n422), .A2(n3147), .B1(n3146), .B2(n3425), .ZN(n2588)
         );
  OAI22_X1 U3396 ( .A1(n422), .A2(n3155), .B1(n3154), .B2(n3425), .ZN(n2596)
         );
  OAI22_X1 U3397 ( .A1(n3576), .A2(n3137), .B1(n3136), .B2(n3425), .ZN(n2578)
         );
  OAI22_X1 U3398 ( .A1(n422), .A2(n3136), .B1(n3135), .B2(n3425), .ZN(n2577)
         );
  OAI22_X1 U3399 ( .A1(n3576), .A2(n3141), .B1(n3140), .B2(n3425), .ZN(n2582)
         );
  OAI22_X1 U3400 ( .A1(n3575), .A2(n3132), .B1(n3131), .B2(n3425), .ZN(n2573)
         );
  NOR2_X1 U3401 ( .A1(n1489), .A2(n1518), .ZN(n3494) );
  NOR2_X1 U3402 ( .A1(n1518), .A2(n1489), .ZN(n788) );
  XNOR2_X2 U3403 ( .A(n1404), .B(n1381), .ZN(n3558) );
  INV_X4 U3404 ( .A(n3676), .ZN(n452) );
  OAI22_X1 U3405 ( .A1(n3603), .A2(n2767), .B1(n3460), .B2(n3280), .ZN(n2197)
         );
  OAI22_X1 U3406 ( .A1(n3602), .A2(n2783), .B1(n2782), .B2(n3460), .ZN(n2213)
         );
  OAI22_X1 U3407 ( .A1(n3602), .A2(n2769), .B1(n2768), .B2(n3459), .ZN(n2199)
         );
  OAI22_X1 U3408 ( .A1(n3602), .A2(n2782), .B1(n2781), .B2(n3459), .ZN(n2212)
         );
  OAI22_X1 U3409 ( .A1(n3602), .A2(n2771), .B1(n2770), .B2(n3460), .ZN(n2201)
         );
  OAI22_X1 U3410 ( .A1(n3602), .A2(n2778), .B1(n2777), .B2(n3460), .ZN(n2208)
         );
  OAI22_X1 U3411 ( .A1(n3603), .A2(n2792), .B1(n2791), .B2(n3460), .ZN(n2222)
         );
  OAI22_X1 U3412 ( .A1(n3602), .A2(n2795), .B1(n2794), .B2(n3459), .ZN(n2225)
         );
  OAI22_X1 U3413 ( .A1(n455), .A2(n2779), .B1(n2778), .B2(n3459), .ZN(n2209)
         );
  OAI22_X1 U3414 ( .A1(n455), .A2(n2784), .B1(n2783), .B2(n3460), .ZN(n2214)
         );
  OAI22_X1 U3415 ( .A1(n455), .A2(n2798), .B1(n2797), .B2(n3459), .ZN(n2228)
         );
  NOR2_X1 U3416 ( .A1(n1612), .A2(n1641), .ZN(n3495) );
  INV_X1 U3417 ( .A(n3730), .ZN(n3496) );
  NOR2_X1 U3418 ( .A1(n1612), .A2(n1641), .ZN(n811) );
  NAND2_X4 U3419 ( .A1(n3583), .A2(n3584), .ZN(n3730) );
  NAND2_X1 U3420 ( .A1(n757), .A2(n760), .ZN(n555) );
  INV_X1 U3421 ( .A(n760), .ZN(n758) );
  OAI21_X1 U3422 ( .B1(n877), .B2(n857), .A(n858), .ZN(n3497) );
  NAND2_X1 U3423 ( .A1(n3498), .A2(n3499), .ZN(n3501) );
  NAND2_X1 U3424 ( .A1(n3500), .A2(n3501), .ZN(n3533) );
  INV_X2 U3425 ( .A(n333), .ZN(n3498) );
  INV_X2 U3426 ( .A(a[10]), .ZN(n3499) );
  XNOR2_X1 U3427 ( .A(n507), .B(n3411), .ZN(n3042) );
  XNOR2_X1 U3428 ( .A(n505), .B(n3411), .ZN(n3043) );
  XNOR2_X1 U3429 ( .A(n503), .B(n3411), .ZN(n3044) );
  XNOR2_X1 U3430 ( .A(n501), .B(n3411), .ZN(n3045) );
  XNOR2_X1 U3431 ( .A(n499), .B(n3411), .ZN(n3046) );
  XNOR2_X1 U3432 ( .A(n497), .B(n3411), .ZN(n3047) );
  XNOR2_X1 U3433 ( .A(n495), .B(n3411), .ZN(n3048) );
  XNOR2_X1 U3434 ( .A(n493), .B(n3411), .ZN(n3049) );
  XNOR2_X1 U3435 ( .A(n491), .B(n3411), .ZN(n3050) );
  XNOR2_X1 U3436 ( .A(n489), .B(n3411), .ZN(n3051) );
  XNOR2_X1 U3437 ( .A(n487), .B(n3411), .ZN(n3052) );
  XNOR2_X1 U3438 ( .A(n485), .B(n3411), .ZN(n3053) );
  XNOR2_X1 U3439 ( .A(n477), .B(n3411), .ZN(n3057) );
  XNOR2_X1 U3440 ( .A(n479), .B(n3411), .ZN(n3056) );
  XNOR2_X1 U3441 ( .A(n483), .B(n3411), .ZN(n3054) );
  XNOR2_X1 U3442 ( .A(n509), .B(n3411), .ZN(n3041) );
  XNOR2_X1 U3443 ( .A(n511), .B(n3411), .ZN(n3040) );
  XNOR2_X1 U3444 ( .A(n513), .B(n3411), .ZN(n3039) );
  XNOR2_X1 U3445 ( .A(n515), .B(n3411), .ZN(n3038) );
  XNOR2_X1 U3446 ( .A(n517), .B(n3411), .ZN(n3037) );
  XNOR2_X1 U3447 ( .A(n519), .B(n3411), .ZN(n3036) );
  XNOR2_X1 U3448 ( .A(n521), .B(n3411), .ZN(n3035) );
  XNOR2_X1 U3449 ( .A(n523), .B(n3411), .ZN(n3034) );
  XNOR2_X1 U3450 ( .A(n525), .B(n3411), .ZN(n3033) );
  XNOR2_X1 U3451 ( .A(n527), .B(n3411), .ZN(n3032) );
  XNOR2_X1 U3452 ( .A(n529), .B(n3411), .ZN(n3031) );
  INV_X1 U3453 ( .A(n3411), .ZN(n3530) );
  OAI22_X1 U3454 ( .A1(n437), .A2(n2976), .B1(n2975), .B2(n387), .ZN(n2412) );
  OAI21_X1 U3455 ( .B1(n800), .B2(n804), .A(n801), .ZN(n799) );
  OAI22_X1 U3456 ( .A1(n3542), .A2(n3084), .B1(n3083), .B2(n3638), .ZN(n2523)
         );
  OAI22_X1 U3457 ( .A1(n3542), .A2(n3079), .B1(n3078), .B2(n3638), .ZN(n2518)
         );
  OR2_X2 U3458 ( .A1(n3737), .A2(n3738), .ZN(n2515) );
  XNOR2_X2 U3459 ( .A(a[16]), .B(n342), .ZN(n3502) );
  OAI22_X1 U3460 ( .A1(n449), .A2(n2863), .B1(n2862), .B2(n399), .ZN(n2295) );
  OAI21_X1 U3461 ( .B1(n3495), .B2(n815), .A(n812), .ZN(n810) );
  NAND2_X1 U3462 ( .A1(n822), .A2(n825), .ZN(n567) );
  INV_X1 U3463 ( .A(n825), .ZN(n823) );
  INV_X4 U3464 ( .A(n3606), .ZN(n3557) );
  AOI21_X1 U3465 ( .B1(n856), .B2(n828), .A(n3444), .ZN(n3503) );
  XOR2_X1 U3466 ( .A(n682), .B(n545), .Z(product[50]) );
  OAI21_X2 U3467 ( .B1(n682), .B2(n680), .A(n681), .ZN(n679) );
  OAI22_X1 U3468 ( .A1(n443), .A2(n2900), .B1(n2899), .B2(n3556), .ZN(n2334)
         );
  OAI22_X1 U3469 ( .A1(n443), .A2(n3284), .B1(n2931), .B2(n3556), .ZN(n2068)
         );
  OAI22_X1 U3470 ( .A1(n443), .A2(n2905), .B1(n2904), .B2(n3556), .ZN(n2339)
         );
  OAI22_X1 U3471 ( .A1(n443), .A2(n2917), .B1(n2916), .B2(n3556), .ZN(n2351)
         );
  OAI22_X1 U3472 ( .A1(n443), .A2(n2912), .B1(n2911), .B2(n3556), .ZN(n2346)
         );
  OAI22_X1 U3473 ( .A1(n443), .A2(n2921), .B1(n2920), .B2(n3556), .ZN(n2355)
         );
  OAI22_X1 U3474 ( .A1(n443), .A2(n2920), .B1(n2919), .B2(n3556), .ZN(n2354)
         );
  OAI22_X1 U3475 ( .A1(n443), .A2(n2923), .B1(n2922), .B2(n3556), .ZN(n2357)
         );
  OAI22_X1 U3476 ( .A1(n443), .A2(n2910), .B1(n2909), .B2(n3556), .ZN(n2344)
         );
  OAI22_X1 U3477 ( .A1(n443), .A2(n2929), .B1(n2928), .B2(n3556), .ZN(n2363)
         );
  OAI22_X1 U3478 ( .A1(n443), .A2(n2926), .B1(n2925), .B2(n3556), .ZN(n2360)
         );
  OAI22_X1 U3479 ( .A1(n443), .A2(n2915), .B1(n2914), .B2(n3556), .ZN(n2349)
         );
  INV_X1 U3480 ( .A(n3604), .ZN(n3605) );
  INV_X1 U3481 ( .A(n3461), .ZN(n796) );
  NOR2_X1 U3482 ( .A1(n777), .A2(n780), .ZN(n3504) );
  NOR2_X2 U3483 ( .A1(n1488), .A2(n3553), .ZN(n780) );
  NOR2_X2 U3484 ( .A1(n811), .A2(n814), .ZN(n809) );
  OAI22_X1 U3485 ( .A1(n449), .A2(n2856), .B1(n2855), .B2(n399), .ZN(n2288) );
  INV_X4 U3486 ( .A(n3672), .ZN(n3541) );
  AOI21_X1 U3487 ( .B1(n3699), .B2(n786), .A(n787), .ZN(n3511) );
  OAI22_X1 U3488 ( .A1(n3649), .A2(n2906), .B1(n2905), .B2(n3556), .ZN(n2340)
         );
  OAI22_X1 U3489 ( .A1(n3649), .A2(n2925), .B1(n2924), .B2(n3556), .ZN(n2359)
         );
  OAI22_X1 U3490 ( .A1(n3649), .A2(n2927), .B1(n2926), .B2(n3556), .ZN(n2361)
         );
  OAI22_X1 U3491 ( .A1(n3649), .A2(n2913), .B1(n2912), .B2(n3556), .ZN(n2347)
         );
  OAI22_X1 U3492 ( .A1(n3649), .A2(n2930), .B1(n2929), .B2(n3556), .ZN(n2364)
         );
  OAI22_X1 U3493 ( .A1(n3649), .A2(n2902), .B1(n2901), .B2(n3556), .ZN(n2336)
         );
  OAI22_X1 U3494 ( .A1(n3649), .A2(n2928), .B1(n2927), .B2(n3556), .ZN(n2362)
         );
  OAI22_X1 U3495 ( .A1(n3649), .A2(n2919), .B1(n2918), .B2(n3556), .ZN(n2353)
         );
  OAI22_X1 U3496 ( .A1(n3649), .A2(n2922), .B1(n2921), .B2(n3556), .ZN(n2356)
         );
  BUF_X1 U3497 ( .A(n3494), .Z(n3505) );
  INV_X4 U3498 ( .A(n3746), .ZN(n3506) );
  AND2_X4 U3499 ( .A1(n3230), .A2(n3453), .ZN(n3746) );
  INV_X4 U3500 ( .A(n3746), .ZN(n458) );
  OAI22_X1 U3501 ( .A1(n3602), .A2(n2774), .B1(n2773), .B2(n3459), .ZN(n2204)
         );
  OAI22_X1 U3502 ( .A1(n3602), .A2(n2775), .B1(n2774), .B2(n3460), .ZN(n2205)
         );
  OAI22_X1 U3503 ( .A1(n3603), .A2(n2791), .B1(n2790), .B2(n3460), .ZN(n2221)
         );
  OAI22_X1 U3504 ( .A1(n3603), .A2(n2790), .B1(n2789), .B2(n3460), .ZN(n2220)
         );
  OAI22_X1 U3505 ( .A1(n3603), .A2(n2780), .B1(n2779), .B2(n3459), .ZN(n2210)
         );
  OAI22_X1 U3506 ( .A1(n3602), .A2(n2787), .B1(n2786), .B2(n3459), .ZN(n2217)
         );
  OAI22_X1 U3507 ( .A1(n3603), .A2(n2777), .B1(n2776), .B2(n3459), .ZN(n2207)
         );
  OAI22_X1 U3508 ( .A1(n3603), .A2(n2788), .B1(n2787), .B2(n3459), .ZN(n2218)
         );
  OAI22_X1 U3509 ( .A1(n455), .A2(n2776), .B1(n2775), .B2(n3459), .ZN(n2206)
         );
  OAI22_X1 U3510 ( .A1(n455), .A2(n2797), .B1(n2796), .B2(n3459), .ZN(n2227)
         );
  OAI22_X1 U3511 ( .A1(n455), .A2(n3280), .B1(n2799), .B2(n3460), .ZN(n2064)
         );
  OAI22_X1 U3512 ( .A1(n3541), .A2(n3091), .B1(n3090), .B2(n3638), .ZN(n2530)
         );
  OAI22_X1 U3513 ( .A1(n3541), .A2(n3069), .B1(n3068), .B2(n3638), .ZN(n2508)
         );
  OAI22_X1 U3514 ( .A1(n3541), .A2(n3075), .B1(n3074), .B2(n3638), .ZN(n2514)
         );
  OAI22_X1 U3515 ( .A1(n3542), .A2(n3094), .B1(n3093), .B2(n3638), .ZN(n2533)
         );
  OAI22_X1 U3516 ( .A1(n3541), .A2(n3088), .B1(n3087), .B2(n3638), .ZN(n2527)
         );
  OAI22_X1 U3517 ( .A1(n3542), .A2(n3086), .B1(n3085), .B2(n3638), .ZN(n2525)
         );
  OAI22_X1 U3518 ( .A1(n3542), .A2(n3095), .B1(n3094), .B2(n3638), .ZN(n2534)
         );
  OAI22_X1 U3519 ( .A1(n3542), .A2(n3632), .B1(n3096), .B2(n3638), .ZN(n2073)
         );
  OAI22_X1 U3520 ( .A1(n3542), .A2(n3071), .B1(n3070), .B2(n3638), .ZN(n2510)
         );
  OAI22_X1 U3521 ( .A1(n3541), .A2(n3074), .B1(n3073), .B2(n3638), .ZN(n2513)
         );
  OAI22_X1 U3522 ( .A1(n3541), .A2(n3067), .B1(n3066), .B2(n3638), .ZN(n2506)
         );
  OAI22_X1 U3523 ( .A1(n3541), .A2(n3083), .B1(n3082), .B2(n3638), .ZN(n2522)
         );
  OAI22_X1 U3524 ( .A1(n3541), .A2(n3087), .B1(n3086), .B2(n3638), .ZN(n2526)
         );
  OAI22_X1 U3525 ( .A1(n3539), .A2(n3121), .B1(n3120), .B2(n375), .ZN(n2561)
         );
  OAI22_X1 U3526 ( .A1(n3539), .A2(n3128), .B1(n3127), .B2(n375), .ZN(n2568)
         );
  OAI22_X1 U3527 ( .A1(n3539), .A2(n3127), .B1(n3126), .B2(n375), .ZN(n2567)
         );
  OAI22_X1 U3528 ( .A1(n3539), .A2(n3126), .B1(n3125), .B2(n375), .ZN(n2566)
         );
  OAI22_X1 U3529 ( .A1(n3539), .A2(n3123), .B1(n3122), .B2(n375), .ZN(n2563)
         );
  OAI22_X1 U3530 ( .A1(n3539), .A2(n3117), .B1(n3116), .B2(n375), .ZN(n2557)
         );
  OAI22_X1 U3531 ( .A1(n3539), .A2(n3112), .B1(n3111), .B2(n375), .ZN(n2552)
         );
  OAI22_X1 U3532 ( .A1(n3539), .A2(n3102), .B1(n3101), .B2(n375), .ZN(n2542)
         );
  OAI22_X1 U3533 ( .A1(n3539), .A2(n3114), .B1(n3113), .B2(n375), .ZN(n2554)
         );
  OAI22_X1 U3534 ( .A1(n3539), .A2(n3103), .B1(n3102), .B2(n375), .ZN(n2543)
         );
  OAI22_X1 U3535 ( .A1(n3539), .A2(n3109), .B1(n3108), .B2(n375), .ZN(n2549)
         );
  OAI22_X1 U3536 ( .A1(n3539), .A2(n3118), .B1(n3117), .B2(n375), .ZN(n2558)
         );
  OAI22_X1 U3537 ( .A1(n3539), .A2(n3113), .B1(n3112), .B2(n375), .ZN(n2553)
         );
  OAI22_X1 U3538 ( .A1(n3539), .A2(n3104), .B1(n3103), .B2(n375), .ZN(n2544)
         );
  NAND2_X1 U3539 ( .A1(n1405), .A2(n1432), .ZN(n3507) );
  NAND2_X1 U3540 ( .A1(n1405), .A2(n1407), .ZN(n3508) );
  NAND2_X1 U3541 ( .A1(n1432), .A2(n1407), .ZN(n3509) );
  NAND3_X1 U3542 ( .A1(n3507), .A2(n3509), .A3(n3508), .ZN(n1402) );
  OAI22_X1 U3543 ( .A1(n3658), .A2(n3060), .B1(n3059), .B2(n381), .ZN(n2498)
         );
  OAI22_X1 U3544 ( .A1(n3658), .A2(n3048), .B1(n3047), .B2(n381), .ZN(n2486)
         );
  OAI22_X1 U3545 ( .A1(n3660), .A2(n3062), .B1(n3061), .B2(n381), .ZN(n2500)
         );
  OAI22_X1 U3546 ( .A1(n3660), .A2(n3042), .B1(n3041), .B2(n381), .ZN(n2480)
         );
  OAI22_X1 U3547 ( .A1(n3660), .A2(n3061), .B1(n3060), .B2(n381), .ZN(n2499)
         );
  OAI22_X1 U3548 ( .A1(n3660), .A2(n3054), .B1(n3053), .B2(n381), .ZN(n2492)
         );
  OAI22_X1 U3549 ( .A1(n3660), .A2(n3059), .B1(n3058), .B2(n381), .ZN(n2497)
         );
  OAI22_X1 U3550 ( .A1(n3660), .A2(n3051), .B1(n3050), .B2(n381), .ZN(n2489)
         );
  OAI22_X1 U3551 ( .A1(n3660), .A2(n3044), .B1(n3043), .B2(n381), .ZN(n2482)
         );
  OAI22_X1 U3552 ( .A1(n3660), .A2(n3052), .B1(n3051), .B2(n381), .ZN(n2490)
         );
  OAI22_X1 U3553 ( .A1(n3659), .A2(n3033), .B1(n3032), .B2(n381), .ZN(n2471)
         );
  OAI22_X1 U3554 ( .A1(n3659), .A2(n3046), .B1(n3045), .B2(n381), .ZN(n2484)
         );
  OAI22_X1 U3555 ( .A1(n3659), .A2(n3053), .B1(n3052), .B2(n381), .ZN(n2491)
         );
  OAI22_X1 U3556 ( .A1(n3660), .A2(n3039), .B1(n3038), .B2(n381), .ZN(n2477)
         );
  OAI22_X1 U3557 ( .A1(n3658), .A2(n3043), .B1(n3042), .B2(n381), .ZN(n2481)
         );
  OAI22_X1 U3558 ( .A1(n3659), .A2(n3041), .B1(n3040), .B2(n381), .ZN(n2479)
         );
  INV_X1 U3559 ( .A(n3607), .ZN(n3510) );
  INV_X4 U3560 ( .A(n3606), .ZN(n3607) );
  OAI21_X1 U3561 ( .B1(n731), .B2(n748), .A(n732), .ZN(n730) );
  NAND2_X2 U3562 ( .A1(n1303), .A2(n1326), .ZN(n748) );
  NOR2_X2 U3563 ( .A1(n1303), .A2(n1326), .ZN(n747) );
  AOI21_X1 U3564 ( .B1(n786), .B2(n799), .A(n787), .ZN(n785) );
  OAI22_X1 U3565 ( .A1(n3575), .A2(n3145), .B1(n3144), .B2(n3425), .ZN(n2586)
         );
  OAI22_X1 U3566 ( .A1(n3576), .A2(n3130), .B1(n3425), .B2(n3615), .ZN(n2571)
         );
  OAI22_X1 U3567 ( .A1(n3576), .A2(n3154), .B1(n3153), .B2(n3425), .ZN(n2595)
         );
  OAI22_X1 U3568 ( .A1(n422), .A2(n3156), .B1(n3155), .B2(n3425), .ZN(n2597)
         );
  OAI22_X1 U3569 ( .A1(n422), .A2(n3159), .B1(n3158), .B2(n3425), .ZN(n2600)
         );
  OAI22_X1 U3570 ( .A1(n3576), .A2(n3161), .B1(n3160), .B2(n3425), .ZN(n2602)
         );
  OAI22_X1 U3571 ( .A1(n422), .A2(n3148), .B1(n3147), .B2(n3425), .ZN(n2589)
         );
  OAI22_X1 U3572 ( .A1(n422), .A2(n3144), .B1(n3143), .B2(n3425), .ZN(n2585)
         );
  OAI22_X1 U3573 ( .A1(n422), .A2(n3139), .B1(n3138), .B2(n3425), .ZN(n2580)
         );
  OAI22_X1 U3574 ( .A1(n3575), .A2(n3133), .B1(n3132), .B2(n3425), .ZN(n2574)
         );
  OAI22_X1 U3575 ( .A1(n3575), .A2(n3143), .B1(n3142), .B2(n3425), .ZN(n2584)
         );
  INV_X4 U3576 ( .A(n3636), .ZN(n3639) );
  NOR2_X2 U3577 ( .A1(n1724), .A2(n1749), .ZN(n834) );
  NAND2_X2 U3578 ( .A1(n3731), .A2(n348), .ZN(n3583) );
  NOR2_X1 U3579 ( .A1(n772), .A2(n769), .ZN(n3512) );
  INV_X1 U3580 ( .A(n3679), .ZN(n3513) );
  NAND2_X2 U3581 ( .A1(n1798), .A2(n1819), .ZN(n850) );
  NOR2_X2 U3582 ( .A1(n1798), .A2(n1819), .ZN(n849) );
  XNOR2_X1 U3583 ( .A(n771), .B(n556), .ZN(product[39]) );
  AOI21_X2 U3584 ( .B1(n783), .B2(n3504), .A(n3705), .ZN(n774) );
  INV_X8 U3585 ( .A(n3690), .ZN(n3666) );
  XOR2_X2 U3586 ( .A(n3514), .B(n2348), .Z(n1577) );
  XOR2_X1 U3587 ( .A(n1571), .B(n1573), .Z(n3515) );
  XOR2_X1 U3588 ( .A(n3515), .B(n1577), .Z(n1563) );
  NAND2_X1 U3589 ( .A1(n2188), .A2(n2124), .ZN(n3516) );
  NAND2_X1 U3590 ( .A1(n2188), .A2(n2348), .ZN(n3517) );
  NAND3_X1 U3591 ( .A1(n3516), .A2(n3517), .A3(n3518), .ZN(n1576) );
  NAND2_X1 U3592 ( .A1(n1571), .A2(n1573), .ZN(n3519) );
  NAND2_X1 U3593 ( .A1(n1571), .A2(n1577), .ZN(n3520) );
  NAND2_X1 U3594 ( .A1(n1573), .A2(n1577), .ZN(n3521) );
  NAND3_X1 U3595 ( .A1(n3519), .A2(n3520), .A3(n3521), .ZN(n1562) );
  OR2_X1 U3596 ( .A1(n2758), .A2(n408), .ZN(n3523) );
  NAND2_X2 U3597 ( .A1(n3522), .A2(n3523), .ZN(n2188) );
  XNOR2_X1 U3598 ( .A(n481), .B(n360), .ZN(n2758) );
  BUF_X4 U3599 ( .A(a[18]), .Z(n3695) );
  INV_X1 U3600 ( .A(n464), .ZN(n3524) );
  INV_X4 U3601 ( .A(n3524), .ZN(n3525) );
  INV_X8 U3602 ( .A(n3744), .ZN(n3526) );
  INV_X1 U3603 ( .A(n3744), .ZN(n414) );
  XNOR2_X1 U3604 ( .A(n701), .B(n3527), .ZN(product[48]) );
  AND2_X1 U3605 ( .A1(n993), .A2(n700), .ZN(n3527) );
  NOR2_X2 U3606 ( .A1(n1431), .A2(n1458), .ZN(n3683) );
  OAI22_X1 U3607 ( .A1(n3477), .A2(n2732), .B1(n2731), .B2(n3607), .ZN(n2160)
         );
  OAI22_X1 U3608 ( .A1(n3477), .A2(n2724), .B1(n2723), .B2(n3607), .ZN(n2152)
         );
  OAI22_X1 U3609 ( .A1(n3477), .A2(n3278), .B1(n2733), .B2(n3607), .ZN(n2062)
         );
  OAI22_X1 U3610 ( .A1(n3476), .A2(n2726), .B1(n2725), .B2(n3607), .ZN(n2154)
         );
  OAI22_X1 U3611 ( .A1(n461), .A2(n2729), .B1(n2728), .B2(n3607), .ZN(n2157)
         );
  OAI22_X1 U3612 ( .A1(n3476), .A2(n2728), .B1(n2727), .B2(n3607), .ZN(n2156)
         );
  OAI22_X1 U3613 ( .A1(n461), .A2(n2722), .B1(n2721), .B2(n3607), .ZN(n2150)
         );
  NOR2_X2 U3614 ( .A1(n3494), .A2(n793), .ZN(n786) );
  OAI22_X1 U3615 ( .A1(n3658), .A2(n3056), .B1(n3055), .B2(n381), .ZN(n2494)
         );
  OAI22_X1 U3616 ( .A1(n3658), .A2(n3036), .B1(n3035), .B2(n381), .ZN(n2474)
         );
  OAI22_X1 U3617 ( .A1(n3660), .A2(n3288), .B1(n3063), .B2(n381), .ZN(n2072)
         );
  OAI22_X1 U3618 ( .A1(n3658), .A2(n3050), .B1(n3049), .B2(n381), .ZN(n2488)
         );
  OAI22_X1 U3619 ( .A1(n3660), .A2(n3058), .B1(n3057), .B2(n381), .ZN(n2496)
         );
  OAI22_X1 U3620 ( .A1(n3658), .A2(n3055), .B1(n3054), .B2(n381), .ZN(n2493)
         );
  OAI22_X1 U3621 ( .A1(n3658), .A2(n3040), .B1(n3039), .B2(n381), .ZN(n2478)
         );
  OAI22_X1 U3622 ( .A1(n3660), .A2(n3057), .B1(n3056), .B2(n381), .ZN(n2495)
         );
  OAI22_X1 U3623 ( .A1(n3658), .A2(n3045), .B1(n3044), .B2(n381), .ZN(n2483)
         );
  OAI22_X1 U3624 ( .A1(n3660), .A2(n3037), .B1(n3036), .B2(n381), .ZN(n2475)
         );
  OAI22_X1 U3625 ( .A1(n3660), .A2(n3032), .B1(n3031), .B2(n381), .ZN(n2470)
         );
  OAI22_X1 U3626 ( .A1(n3660), .A2(n3049), .B1(n3048), .B2(n381), .ZN(n2487)
         );
  OAI22_X1 U3627 ( .A1(n3660), .A2(n3034), .B1(n3033), .B2(n381), .ZN(n2472)
         );
  OAI22_X1 U3628 ( .A1(n3660), .A2(n3031), .B1(n381), .B2(n3288), .ZN(n2469)
         );
  OAI22_X1 U3629 ( .A1(n3660), .A2(n3035), .B1(n3034), .B2(n381), .ZN(n2473)
         );
  OAI22_X1 U3630 ( .A1(n3660), .A2(n3038), .B1(n3037), .B2(n381), .ZN(n2476)
         );
  OAI22_X1 U3631 ( .A1(n446), .A2(n3283), .B1(n2898), .B2(n396), .ZN(n2067) );
  OAI22_X1 U3632 ( .A1(n446), .A2(n2881), .B1(n2880), .B2(n396), .ZN(n2314) );
  OAI22_X1 U3633 ( .A1(n446), .A2(n2879), .B1(n2878), .B2(n396), .ZN(n2312) );
  OAI22_X1 U3634 ( .A1(n446), .A2(n2887), .B1(n2886), .B2(n396), .ZN(n2320) );
  OAI22_X1 U3635 ( .A1(n446), .A2(n2882), .B1(n2881), .B2(n396), .ZN(n2315) );
  OAI22_X1 U3636 ( .A1(n446), .A2(n2877), .B1(n2876), .B2(n396), .ZN(n2310) );
  OAI22_X1 U3637 ( .A1(n446), .A2(n2888), .B1(n2887), .B2(n396), .ZN(n2321) );
  OAI22_X1 U3638 ( .A1(n446), .A2(n2896), .B1(n2895), .B2(n396), .ZN(n2329) );
  OAI21_X1 U3639 ( .B1(n3683), .B2(n781), .A(n778), .ZN(n3528) );
  NAND2_X2 U3640 ( .A1(n1459), .A2(n1488), .ZN(n781) );
  NOR2_X1 U3641 ( .A1(n727), .A2(n613), .ZN(n611) );
  OR2_X4 U3642 ( .A1(n3529), .A2(a[0]), .ZN(n419) );
  XNOR2_X2 U3643 ( .A(a[0]), .B(n321), .ZN(n3529) );
  XOR2_X2 U3644 ( .A(n3750), .B(n3577), .Z(n3749) );
  INV_X1 U3645 ( .A(n419), .ZN(n3754) );
  NAND2_X1 U3646 ( .A1(a[30]), .A2(n3645), .ZN(n3646) );
  INV_X2 U3647 ( .A(n363), .ZN(n3645) );
  INV_X4 U3648 ( .A(a[26]), .ZN(n3635) );
  OAI22_X1 U3649 ( .A1(n3680), .A2(n3016), .B1(n3015), .B2(n384), .ZN(n2453)
         );
  OAI22_X1 U3650 ( .A1(n3680), .A2(n2999), .B1(n2998), .B2(n384), .ZN(n2436)
         );
  OAI22_X1 U3651 ( .A1(n3680), .A2(n3029), .B1(n3028), .B2(n384), .ZN(n2466)
         );
  OAI22_X1 U3652 ( .A1(n3680), .A2(n3287), .B1(n3030), .B2(n384), .ZN(n2071)
         );
  OAI22_X1 U3653 ( .A1(n3680), .A2(n3011), .B1(n3010), .B2(n384), .ZN(n2448)
         );
  OAI22_X1 U3654 ( .A1(n3680), .A2(n3010), .B1(n3009), .B2(n384), .ZN(n2447)
         );
  OAI22_X1 U3655 ( .A1(n3680), .A2(n3023), .B1(n3022), .B2(n384), .ZN(n2460)
         );
  OAI22_X1 U3656 ( .A1(n3680), .A2(n3000), .B1(n2999), .B2(n384), .ZN(n2437)
         );
  OAI22_X1 U3657 ( .A1(n3680), .A2(n3024), .B1(n3023), .B2(n384), .ZN(n2461)
         );
  OAI22_X1 U3658 ( .A1(n3680), .A2(n3027), .B1(n3026), .B2(n384), .ZN(n2464)
         );
  OAI22_X1 U3659 ( .A1(n3680), .A2(n3003), .B1(n3002), .B2(n384), .ZN(n2440)
         );
  OAI22_X1 U3660 ( .A1(n3680), .A2(n3028), .B1(n3027), .B2(n384), .ZN(n2465)
         );
  OAI22_X1 U3661 ( .A1(n3680), .A2(n3008), .B1(n3007), .B2(n384), .ZN(n2445)
         );
  OAI22_X1 U3662 ( .A1(n3680), .A2(n3020), .B1(n3019), .B2(n384), .ZN(n2457)
         );
  OAI22_X1 U3663 ( .A1(n3680), .A2(n3025), .B1(n3024), .B2(n384), .ZN(n2462)
         );
  OAI22_X1 U3664 ( .A1(n3680), .A2(n3007), .B1(n3006), .B2(n384), .ZN(n2444)
         );
  OAI22_X1 U3665 ( .A1(n3680), .A2(n3026), .B1(n3025), .B2(n384), .ZN(n2463)
         );
  AND2_X2 U3666 ( .A1(n3543), .A2(n3544), .ZN(n766) );
  OAI21_X2 U3667 ( .B1(n3653), .B2(n688), .A(n689), .ZN(n687) );
  AOI21_X2 U3668 ( .B1(n687), .B2(n673), .A(n676), .ZN(n672) );
  INV_X4 U3669 ( .A(a[28]), .ZN(n3656) );
  OAI22_X1 U3670 ( .A1(n464), .A2(n2697), .B1(n2696), .B2(n3526), .ZN(n2124)
         );
  XOR2_X2 U3671 ( .A(n3729), .B(n3604), .Z(n3728) );
  OAI21_X1 U3672 ( .B1(n3503), .B2(n807), .A(n808), .ZN(n3532) );
  OAI21_X1 U3673 ( .B1(n3443), .B2(n807), .A(n808), .ZN(n3618) );
  NAND2_X1 U3674 ( .A1(n3678), .A2(n672), .ZN(n670) );
  OAI22_X1 U3675 ( .A1(n464), .A2(n2693), .B1(n2692), .B2(n3526), .ZN(n2120)
         );
  NAND2_X1 U3676 ( .A1(n3678), .A2(n672), .ZN(n3621) );
  INV_X1 U3677 ( .A(n3725), .ZN(n411) );
  INV_X8 U3678 ( .A(n3622), .ZN(n3535) );
  INV_X1 U3679 ( .A(n3742), .ZN(n3536) );
  OAI21_X1 U3680 ( .B1(n3511), .B2(n765), .A(n766), .ZN(n764) );
  INV_X1 U3681 ( .A(n3448), .ZN(n3537) );
  INV_X4 U3682 ( .A(n3448), .ZN(n3539) );
  INV_X4 U3683 ( .A(n3448), .ZN(n3538) );
  INV_X1 U3684 ( .A(n3686), .ZN(n3540) );
  INV_X8 U3685 ( .A(n3686), .ZN(n387) );
  NAND2_X1 U3686 ( .A1(a[12]), .A2(n3641), .ZN(n3642) );
  OAI22_X1 U3687 ( .A1(n3542), .A2(n3065), .B1(n3064), .B2(n3639), .ZN(n2504)
         );
  OAI22_X1 U3688 ( .A1(n3542), .A2(n3081), .B1(n3080), .B2(n3638), .ZN(n2520)
         );
  OAI22_X1 U3689 ( .A1(n3542), .A2(n3073), .B1(n3072), .B2(n3639), .ZN(n2512)
         );
  OAI22_X1 U3690 ( .A1(n3542), .A2(n3078), .B1(n3077), .B2(n3638), .ZN(n2517)
         );
  INV_X4 U3691 ( .A(n3672), .ZN(n3542) );
  INV_X1 U3692 ( .A(n3672), .ZN(n428) );
  AND2_X4 U3693 ( .A1(n3240), .A2(n3637), .ZN(n3672) );
  OAI22_X1 U3694 ( .A1(n434), .A2(n3004), .B1(n3003), .B2(n384), .ZN(n2441) );
  OAI22_X1 U3695 ( .A1(n434), .A2(n3014), .B1(n3013), .B2(n384), .ZN(n2451) );
  OAI22_X1 U3696 ( .A1(n434), .A2(n3015), .B1(n3014), .B2(n384), .ZN(n2452) );
  OAI22_X1 U3697 ( .A1(n434), .A2(n3013), .B1(n3012), .B2(n384), .ZN(n2450) );
  OAI22_X1 U3698 ( .A1(n434), .A2(n3001), .B1(n3000), .B2(n384), .ZN(n2438) );
  OAI22_X1 U3699 ( .A1(n434), .A2(n3002), .B1(n3001), .B2(n384), .ZN(n2439) );
  OAI22_X1 U3700 ( .A1(n434), .A2(n2998), .B1(n384), .B2(n3287), .ZN(n2435) );
  OAI22_X1 U3701 ( .A1(n434), .A2(n3009), .B1(n3008), .B2(n384), .ZN(n2446) );
  OAI22_X1 U3702 ( .A1(n434), .A2(n3021), .B1(n3020), .B2(n384), .ZN(n2458) );
  OAI22_X1 U3703 ( .A1(n434), .A2(n3022), .B1(n3021), .B2(n384), .ZN(n2459) );
  OAI22_X1 U3704 ( .A1(n434), .A2(n3017), .B1(n3016), .B2(n384), .ZN(n2454) );
  OAI22_X1 U3705 ( .A1(n434), .A2(n3018), .B1(n3017), .B2(n384), .ZN(n2455) );
  OAI22_X1 U3706 ( .A1(n434), .A2(n3019), .B1(n3018), .B2(n384), .ZN(n2456) );
  NAND2_X1 U3707 ( .A1(n3528), .A2(n3512), .ZN(n3543) );
  INV_X1 U3708 ( .A(n768), .ZN(n3544) );
  AOI21_X1 U3709 ( .B1(n670), .B2(n654), .A(n655), .ZN(n3546) );
  AOI21_X1 U3710 ( .B1(n3621), .B2(n654), .A(n655), .ZN(n3545) );
  AOI21_X1 U3711 ( .B1(n670), .B2(n654), .A(n655), .ZN(n653) );
  XOR2_X1 U3712 ( .A(n1671), .B(n1646), .Z(n3547) );
  NAND2_X1 U3713 ( .A1(n1644), .A2(n1671), .ZN(n3548) );
  NAND2_X1 U3714 ( .A1(n1644), .A2(n1646), .ZN(n3549) );
  NAND2_X1 U3715 ( .A1(n1671), .A2(n1646), .ZN(n3550) );
  NAND3_X1 U3716 ( .A1(n3548), .A2(n3550), .A3(n3549), .ZN(n1641) );
  AOI21_X1 U3717 ( .B1(n999), .B2(n749), .A(n746), .ZN(n3551) );
  OAI21_X2 U3718 ( .B1(n3665), .B2(n750), .A(n751), .ZN(n749) );
  AOI21_X1 U3719 ( .B1(n749), .B2(n999), .A(n746), .ZN(n744) );
  XNOR2_X1 U3720 ( .A(n1492), .B(n3552), .ZN(n1461) );
  XNOR2_X1 U3721 ( .A(n1494), .B(n1465), .ZN(n3552) );
  INV_X4 U3722 ( .A(n3502), .ZN(n3554) );
  INV_X2 U3723 ( .A(n3554), .ZN(n3555) );
  FA_X1 U3724 ( .A(n1490), .B(n1463), .CI(n1461), .S(n3553) );
  INV_X4 U3725 ( .A(n3690), .ZN(n446) );
  OR2_X2 U3726 ( .A1(n3697), .A2(n3696), .ZN(n2516) );
  XNOR2_X1 U3727 ( .A(n698), .B(n546), .ZN(product[49]) );
  INV_X8 U3728 ( .A(n3554), .ZN(n3556) );
  AND2_X2 U3729 ( .A1(n3600), .A2(n3601), .ZN(n808) );
  NAND2_X2 U3730 ( .A1(n3642), .A2(n3643), .ZN(n3686) );
  XNOR2_X2 U3731 ( .A(n1379), .B(n3558), .ZN(n1377) );
  NOR2_X1 U3732 ( .A1(n777), .A2(n780), .ZN(n775) );
  NAND2_X1 U3733 ( .A1(n995), .A2(n716), .ZN(n549) );
  AOI21_X2 U3734 ( .B1(n995), .B2(n721), .A(n714), .ZN(n712) );
  NAND2_X2 U3735 ( .A1(n996), .A2(n995), .ZN(n711) );
  NAND2_X1 U3736 ( .A1(n1219), .A2(n1238), .ZN(n716) );
  NOR2_X1 U3737 ( .A1(n1219), .A2(n1238), .ZN(n715) );
  NAND2_X1 U3738 ( .A1(n753), .A2(n3475), .ZN(n3559) );
  AND2_X2 U3739 ( .A1(n3559), .A2(n3442), .ZN(n3653) );
  BUF_X1 U3740 ( .A(n772), .Z(n3560) );
  INV_X1 U3741 ( .A(n3709), .ZN(n3561) );
  INV_X8 U3742 ( .A(n3652), .ZN(n402) );
  NAND2_X1 U3743 ( .A1(n1492), .A2(n1494), .ZN(n3562) );
  NAND2_X1 U3744 ( .A1(n1492), .A2(n1465), .ZN(n3563) );
  NAND2_X1 U3745 ( .A1(n1494), .A2(n1465), .ZN(n3564) );
  NAND3_X2 U3746 ( .A1(n3562), .A2(n3564), .A3(n3563), .ZN(n1460) );
  INV_X1 U3747 ( .A(n3445), .ZN(n1000) );
  NAND2_X1 U3748 ( .A1(n1327), .A2(n1350), .ZN(n755) );
  OAI21_X1 U3749 ( .B1(n3758), .B2(n3745), .A(n3712), .ZN(n2332) );
  NAND2_X1 U3750 ( .A1(n1379), .A2(n1404), .ZN(n3565) );
  NAND2_X1 U3751 ( .A1(n1379), .A2(n1381), .ZN(n3566) );
  NAND2_X1 U3752 ( .A1(n1404), .A2(n1381), .ZN(n3567) );
  NAND3_X1 U3753 ( .A1(n3565), .A2(n3567), .A3(n3566), .ZN(n1376) );
  NAND2_X2 U3754 ( .A1(n1351), .A2(n1376), .ZN(n760) );
  NAND2_X1 U3755 ( .A1(n690), .A2(n615), .ZN(n613) );
  INV_X2 U3756 ( .A(n3651), .ZN(n3652) );
  BUF_X1 U3757 ( .A(n803), .Z(n3569) );
  NAND2_X1 U3758 ( .A1(n3743), .A2(n339), .ZN(n3572) );
  NAND2_X1 U3759 ( .A1(n3570), .A2(n3571), .ZN(n3573) );
  NAND2_X1 U3760 ( .A1(n3572), .A2(n3573), .ZN(n3742) );
  INV_X1 U3761 ( .A(n3743), .ZN(n3570) );
  NOR2_X1 U3762 ( .A1(n1582), .A2(n1611), .ZN(n803) );
  INV_X4 U3763 ( .A(a[14]), .ZN(n3743) );
  INV_X1 U3764 ( .A(n3742), .ZN(n3608) );
  INV_X1 U3765 ( .A(n3569), .ZN(n1009) );
  XNOR2_X1 U3766 ( .A(n2539), .B(n3574), .ZN(n1545) );
  XNOR2_X1 U3767 ( .A(n2155), .B(n2123), .ZN(n3574) );
  NAND2_X4 U3768 ( .A1(n3242), .A2(n372), .ZN(n3576) );
  INV_X2 U3769 ( .A(n3577), .ZN(n3578) );
  BUF_X1 U3770 ( .A(n3497), .Z(n3579) );
  OAI21_X2 U3771 ( .B1(n805), .B2(n784), .A(n3619), .ZN(n783) );
  XNOR2_X1 U3772 ( .A(n1462), .B(n3580), .ZN(n1433) );
  XNOR2_X1 U3773 ( .A(n1437), .B(n1464), .ZN(n3580) );
  NAND2_X1 U3774 ( .A1(n3581), .A2(n3582), .ZN(n3584) );
  INV_X1 U3775 ( .A(n3409), .ZN(n3581) );
  INV_X1 U3776 ( .A(n348), .ZN(n3582) );
  NAND2_X2 U3777 ( .A1(n3655), .A2(n997), .ZN(n731) );
  BUF_X1 U3778 ( .A(n773), .Z(n3585) );
  NAND2_X1 U3779 ( .A1(n345), .A2(n3587), .ZN(n3588) );
  NAND2_X1 U3780 ( .A1(n3586), .A2(a[18]), .ZN(n3589) );
  NAND2_X1 U3781 ( .A1(n3588), .A2(n3589), .ZN(n3679) );
  INV_X2 U3782 ( .A(n345), .ZN(n3586) );
  BUF_X4 U3783 ( .A(n345), .Z(n3712) );
  XNOR2_X1 U3784 ( .A(n497), .B(n345), .ZN(n2915) );
  XNOR2_X1 U3785 ( .A(n477), .B(n345), .ZN(n2925) );
  XOR2_X1 U3786 ( .A(n2607), .B(n2127), .Z(n3590) );
  XOR2_X1 U3787 ( .A(n2159), .B(n3590), .Z(n1668) );
  NAND2_X1 U3788 ( .A1(n2159), .A2(n3447), .ZN(n3591) );
  NAND2_X1 U3789 ( .A1(n2159), .A2(n2127), .ZN(n3592) );
  NAND2_X1 U3790 ( .A1(n3447), .A2(n2127), .ZN(n3593) );
  NAND3_X1 U3791 ( .A1(n3591), .A2(n3593), .A3(n3592), .ZN(n1667) );
  OR2_X2 U3792 ( .A1(n3476), .A2(n2731), .ZN(n3594) );
  OR2_X1 U3793 ( .A1(n2730), .A2(n3607), .ZN(n3595) );
  NAND2_X2 U3794 ( .A1(n3594), .A2(n3595), .ZN(n2159) );
  OAI22_X1 U3795 ( .A1(n419), .A2(n3165), .B1(n3164), .B2(n369), .ZN(n2607) );
  NOR2_X1 U3796 ( .A1(n3526), .A2(n3440), .ZN(n2127) );
  XNOR2_X1 U3797 ( .A(n471), .B(n363), .ZN(n2730) );
  NAND2_X1 U3798 ( .A1(n3596), .A2(n3597), .ZN(n3599) );
  INV_X1 U3799 ( .A(n3635), .ZN(n3596) );
  INV_X1 U3800 ( .A(n357), .ZN(n3597) );
  NAND2_X1 U3801 ( .A1(n818), .A2(n809), .ZN(n3600) );
  INV_X1 U3802 ( .A(n810), .ZN(n3601) );
  INV_X4 U3803 ( .A(n354), .ZN(n3604) );
  INV_X2 U3804 ( .A(n411), .ZN(n3606) );
  NAND2_X1 U3805 ( .A1(n1008), .A2(n801), .ZN(n562) );
  OAI22_X1 U3806 ( .A1(n449), .A2(n2846), .B1(n2845), .B2(n399), .ZN(n2278) );
  OAI21_X1 U3807 ( .B1(n3755), .B2(n3749), .A(n324), .ZN(n2570) );
  INV_X2 U3808 ( .A(n3608), .ZN(n3609) );
  NAND2_X1 U3809 ( .A1(a[22]), .A2(n3611), .ZN(n3612) );
  NAND2_X1 U3810 ( .A1(n3610), .A2(n351), .ZN(n3613) );
  NAND2_X1 U3811 ( .A1(n3612), .A2(n3613), .ZN(n3709) );
  OAI21_X2 U3812 ( .B1(n665), .B2(n663), .A(n664), .ZN(n662) );
  NAND2_X1 U3813 ( .A1(n3614), .A2(n3615), .ZN(n3617) );
  NAND2_X2 U3814 ( .A1(n3616), .A2(n3617), .ZN(n3747) );
  INV_X1 U3815 ( .A(n3748), .ZN(n3614) );
  INV_X1 U3816 ( .A(n324), .ZN(n3615) );
  OAI21_X1 U3817 ( .B1(n827), .B2(n807), .A(n808), .ZN(n806) );
  OAI22_X1 U3818 ( .A1(n449), .A2(n2848), .B1(n2847), .B2(n399), .ZN(n2280) );
  BUF_X1 U3819 ( .A(n3511), .Z(n3619) );
  XNOR2_X1 U3820 ( .A(n595), .B(n3620), .ZN(product[63]) );
  XNOR2_X1 U3821 ( .A(n1042), .B(n1041), .ZN(n3620) );
  XNOR2_X1 U3822 ( .A(n662), .B(n541), .ZN(product[54]) );
  INV_X1 U3823 ( .A(n422), .ZN(n3755) );
  OAI22_X1 U3824 ( .A1(n3575), .A2(n3135), .B1(n3134), .B2(n3425), .ZN(n2576)
         );
  OAI21_X1 U3825 ( .B1(n3759), .B2(n3728), .A(n357), .ZN(n2196) );
  INV_X8 U3826 ( .A(n3730), .ZN(n399) );
  OAI22_X1 U3827 ( .A1(n434), .A2(n3006), .B1(n3005), .B2(n384), .ZN(n2443) );
  INV_X8 U3828 ( .A(n3622), .ZN(n440) );
  OAI22_X1 U3829 ( .A1(n3537), .A2(n3097), .B1(n375), .B2(n3290), .ZN(n2537)
         );
  OAI21_X1 U3830 ( .B1(n855), .B2(n842), .A(n3434), .ZN(n841) );
  NAND2_X1 U3831 ( .A1(n1489), .A2(n1518), .ZN(n789) );
  XNOR2_X1 U3832 ( .A(n1491), .B(n3704), .ZN(n1489) );
  NAND2_X1 U3833 ( .A1(n2539), .A2(n2155), .ZN(n3623) );
  NAND2_X1 U3834 ( .A1(n2539), .A2(n2123), .ZN(n3624) );
  NAND2_X1 U3835 ( .A1(n2155), .A2(n2123), .ZN(n3625) );
  NAND3_X1 U3836 ( .A1(n3623), .A2(n3625), .A3(n3624), .ZN(n1544) );
  OR2_X1 U3837 ( .A1(n3539), .A2(n3099), .ZN(n3626) );
  OR2_X1 U3838 ( .A1(n3098), .A2(n375), .ZN(n3627) );
  NAND2_X1 U3839 ( .A1(n3626), .A2(n3627), .ZN(n2539) );
  OAI22_X1 U3840 ( .A1(n464), .A2(n2696), .B1(n2695), .B2(n3526), .ZN(n2123)
         );
  OAI22_X1 U3841 ( .A1(n3476), .A2(n2727), .B1(n2726), .B2(n3557), .ZN(n2155)
         );
  XNOR2_X1 U3842 ( .A(n525), .B(n3482), .ZN(n3099) );
  XNOR2_X1 U3843 ( .A(n527), .B(n3726), .ZN(n3098) );
  INV_X2 U3844 ( .A(n3667), .ZN(n3668) );
  OR2_X2 U3845 ( .A1(n3733), .A2(n3734), .ZN(n2313) );
  INV_X8 U3846 ( .A(n3668), .ZN(n396) );
  OAI21_X1 U3847 ( .B1(n788), .B2(n794), .A(n789), .ZN(n787) );
  NAND2_X1 U3848 ( .A1(n859), .A2(n867), .ZN(n857) );
  NAND2_X1 U3849 ( .A1(n1462), .A2(n1437), .ZN(n3628) );
  NAND2_X1 U3850 ( .A1(n1462), .A2(n1464), .ZN(n3629) );
  NAND2_X1 U3851 ( .A1(n1437), .A2(n1464), .ZN(n3630) );
  NAND3_X1 U3852 ( .A1(n3628), .A2(n3630), .A3(n3629), .ZN(n1432) );
  NAND2_X2 U3853 ( .A1(n3752), .A2(n330), .ZN(n3633) );
  NAND2_X1 U3854 ( .A1(n3631), .A2(n3632), .ZN(n3634) );
  INV_X1 U3855 ( .A(n3752), .ZN(n3631) );
  INV_X8 U3856 ( .A(n3687), .ZN(n408) );
  INV_X1 U3857 ( .A(n3691), .ZN(n3637) );
  INV_X4 U3858 ( .A(n3636), .ZN(n3638) );
  NAND2_X2 U3859 ( .A1(n3644), .A2(n363), .ZN(n3647) );
  NAND2_X2 U3860 ( .A1(n3646), .A2(n3647), .ZN(n3744) );
  OAI22_X1 U3861 ( .A1(n3671), .A2(n2819), .B1(n2818), .B2(n402), .ZN(n2250)
         );
  OAI22_X1 U3862 ( .A1(n452), .A2(n2815), .B1(n2814), .B2(n402), .ZN(n2246) );
  OAI22_X1 U3863 ( .A1(n452), .A2(n2828), .B1(n2827), .B2(n402), .ZN(n2259) );
  OAI22_X1 U3864 ( .A1(n452), .A2(n2829), .B1(n2828), .B2(n402), .ZN(n2260) );
  OAI22_X1 U3865 ( .A1(n3671), .A2(n2820), .B1(n2819), .B2(n402), .ZN(n2251)
         );
  OAI22_X1 U3866 ( .A1(n3671), .A2(n2821), .B1(n2820), .B2(n402), .ZN(n2252)
         );
  OAI22_X1 U3867 ( .A1(n452), .A2(n2825), .B1(n2824), .B2(n402), .ZN(n2256) );
  OAI22_X1 U3868 ( .A1(n3671), .A2(n2811), .B1(n2810), .B2(n402), .ZN(n2242)
         );
  OAI22_X1 U3869 ( .A1(n3671), .A2(n2824), .B1(n2823), .B2(n402), .ZN(n2255)
         );
  OAI22_X1 U3870 ( .A1(n3671), .A2(n2822), .B1(n2821), .B2(n402), .ZN(n2253)
         );
  OAI22_X1 U3871 ( .A1(n3671), .A2(n2823), .B1(n2822), .B2(n402), .ZN(n2254)
         );
  OAI22_X1 U3872 ( .A1(n3671), .A2(n2826), .B1(n2825), .B2(n402), .ZN(n2257)
         );
  OAI22_X1 U3873 ( .A1(n3671), .A2(n2817), .B1(n2816), .B2(n402), .ZN(n2248)
         );
  OAI22_X1 U3874 ( .A1(n3671), .A2(n2805), .B1(n2804), .B2(n402), .ZN(n2236)
         );
  OAI22_X1 U3875 ( .A1(n452), .A2(n2830), .B1(n2829), .B2(n402), .ZN(n2261) );
  BUF_X1 U3876 ( .A(n3443), .Z(n3727) );
  OAI21_X1 U3877 ( .B1(n3661), .B2(n3730), .A(n351), .ZN(n2264) );
  OAI22_X1 U3878 ( .A1(n3436), .A2(n2989), .B1(n2988), .B2(n387), .ZN(n2425)
         );
  INV_X8 U3879 ( .A(n3747), .ZN(n375) );
  AOI21_X1 U3880 ( .B1(n603), .B2(n980), .A(n600), .ZN(n3648) );
  NAND2_X4 U3881 ( .A1(n3235), .A2(n3555), .ZN(n3650) );
  NAND2_X4 U3882 ( .A1(n3235), .A2(n3555), .ZN(n3649) );
  AOI21_X1 U3883 ( .B1(n603), .B2(n980), .A(n600), .ZN(n598) );
  INV_X1 U3884 ( .A(n3709), .ZN(n3651) );
  AOI21_X1 U3885 ( .B1(n753), .B2(n3475), .A(n730), .ZN(n728) );
  INV_X1 U3886 ( .A(n686), .ZN(n684) );
  OR2_X4 U3887 ( .A1(n1281), .A2(n1302), .ZN(n3655) );
  INV_X4 U3888 ( .A(n3655), .ZN(n738) );
  XNOR2_X2 U3889 ( .A(n1521), .B(n3657), .ZN(n1519) );
  XNOR2_X2 U3890 ( .A(n1552), .B(n1523), .ZN(n3657) );
  INV_X1 U3891 ( .A(n3462), .ZN(n3658) );
  INV_X4 U3892 ( .A(n3462), .ZN(n3660) );
  OAI22_X1 U3893 ( .A1(n3659), .A2(n3047), .B1(n3046), .B2(n381), .ZN(n2485)
         );
  INV_X1 U3894 ( .A(n3660), .ZN(n3757) );
  OAI21_X1 U3895 ( .B1(n3756), .B2(n3747), .A(n3740), .ZN(n2536) );
  INV_X1 U3896 ( .A(n834), .ZN(n832) );
  INV_X1 U3897 ( .A(n800), .ZN(n1008) );
  NOR2_X2 U3898 ( .A1(n803), .A2(n800), .ZN(n798) );
  AOI21_X2 U3899 ( .B1(n997), .B2(n741), .A(n734), .ZN(n732) );
  INV_X1 U3900 ( .A(n739), .ZN(n741) );
  AOI21_X2 U3901 ( .B1(n691), .B2(n615), .A(n616), .ZN(n614) );
  INV_X1 U3902 ( .A(n687), .ZN(n685) );
  AND2_X2 U3903 ( .A1(n3233), .A2(n3496), .ZN(n3661) );
  INV_X8 U3904 ( .A(n3661), .ZN(n449) );
  INV_X8 U3905 ( .A(n3609), .ZN(n390) );
  AOI21_X2 U3906 ( .B1(n3618), .B2(n763), .A(n3534), .ZN(n3670) );
  NOR2_X2 U3907 ( .A1(n727), .A2(n688), .ZN(n686) );
  OAI22_X1 U3908 ( .A1(n437), .A2(n2970), .B1(n2969), .B2(n387), .ZN(n2406) );
  NAND2_X1 U3909 ( .A1(n1551), .A2(n1581), .ZN(n801) );
  XOR2_X1 U3910 ( .A(n805), .B(n563), .Z(product[32]) );
  OAI21_X1 U3911 ( .B1(n805), .B2(n796), .A(n797), .ZN(n795) );
  OAI21_X1 U3912 ( .B1(n3757), .B2(n3751), .A(n3531), .ZN(n2468) );
  NAND2_X1 U3913 ( .A1(n997), .A2(n736), .ZN(n551) );
  NAND2_X1 U3914 ( .A1(n1259), .A2(n1280), .ZN(n736) );
  NOR2_X1 U3915 ( .A1(n1259), .A2(n1280), .ZN(n735) );
  OR2_X2 U3916 ( .A1(n3707), .A2(n3708), .ZN(n2507) );
  INV_X1 U3917 ( .A(n3654), .ZN(n726) );
  NAND2_X1 U3918 ( .A1(n1521), .A2(n1552), .ZN(n3662) );
  NAND2_X1 U3919 ( .A1(n1521), .A2(n1523), .ZN(n3663) );
  NAND2_X1 U3920 ( .A1(n1552), .A2(n1523), .ZN(n3664) );
  NAND3_X1 U3921 ( .A1(n3662), .A2(n3664), .A3(n3663), .ZN(n1518) );
  AOI21_X1 U3922 ( .B1(n3532), .B2(n763), .A(n3534), .ZN(n3665) );
  INV_X1 U3923 ( .A(n3679), .ZN(n3667) );
  NOR2_X1 U3924 ( .A1(n1377), .A2(n1402), .ZN(n3669) );
  AOI21_X1 U3925 ( .B1(n806), .B2(n763), .A(n764), .ZN(n531) );
  AND2_X2 U3926 ( .A1(n3228), .A2(n414), .ZN(n3673) );
  INV_X8 U3927 ( .A(n3673), .ZN(n464) );
  OAI21_X1 U3928 ( .B1(n3622), .B2(n3609), .A(n342), .ZN(n2366) );
  XNOR2_X1 U3929 ( .A(n1759), .B(n3675), .ZN(n1730) );
  XNOR2_X1 U3930 ( .A(n1736), .B(n1738), .ZN(n3675) );
  OAI21_X1 U3931 ( .B1(n3690), .B2(n3668), .A(n348), .ZN(n2298) );
  OAI22_X1 U3932 ( .A1(n458), .A2(n2763), .B1(n2762), .B2(n408), .ZN(n2192) );
  OAI21_X1 U3933 ( .B1(n3724), .B2(n3686), .A(n339), .ZN(n2400) );
  INV_X1 U3934 ( .A(n3532), .ZN(n805) );
  XNOR2_X2 U3935 ( .A(n1553), .B(n3677), .ZN(n1551) );
  XNOR2_X1 U3936 ( .A(n1583), .B(n1555), .ZN(n3677) );
  OAI21_X1 U3937 ( .B1(n3673), .B2(n3744), .A(n3410), .ZN(n3760) );
  OAI21_X1 U3938 ( .B1(n3676), .B2(n3652), .A(n3605), .ZN(n2230) );
  NAND2_X1 U3939 ( .A1(n3698), .A2(n770), .ZN(n556) );
  OAI21_X1 U3940 ( .B1(n3746), .B2(n3687), .A(n360), .ZN(n2162) );
  NAND2_X1 U3941 ( .A1(n1724), .A2(n1749), .ZN(n835) );
  OAI21_X1 U3942 ( .B1(n3674), .B2(n3510), .A(n363), .ZN(n2128) );
  OAI21_X1 U3943 ( .B1(n805), .B2(n3569), .A(n804), .ZN(n802) );
  NAND2_X1 U3944 ( .A1(n1009), .A2(n804), .ZN(n563) );
  NAND2_X1 U3945 ( .A1(n611), .A2(n981), .ZN(n604) );
  NOR2_X1 U3946 ( .A1(n2662), .A2(n3455), .ZN(n1428) );
  INV_X1 U3947 ( .A(n1428), .ZN(n1429) );
  OR2_X2 U3948 ( .A1(n531), .A2(n671), .ZN(n3678) );
  OAI21_X1 U3949 ( .B1(n3665), .B2(n604), .A(n605), .ZN(n603) );
  INV_X16 U3950 ( .A(a[0]), .ZN(n369) );
  INV_X4 U3951 ( .A(n3741), .ZN(n3680) );
  INV_X1 U3952 ( .A(n907), .ZN(n1026) );
  OAI21_X2 U3953 ( .B1(n907), .B2(n913), .A(n908), .ZN(n906) );
  NAND2_X1 U3954 ( .A1(n1964), .A2(n1977), .ZN(n908) );
  NAND2_X1 U3955 ( .A1(n1003), .A2(n3585), .ZN(n557) );
  NAND2_X1 U3956 ( .A1(n1403), .A2(n1430), .ZN(n773) );
  AOI21_X1 U3957 ( .B1(n817), .B2(n826), .A(n3446), .ZN(n816) );
  NOR2_X1 U3958 ( .A1(n819), .A2(n824), .ZN(n817) );
  FA_X1 U3959 ( .A(n1460), .B(n1435), .CI(n1433), .S(n3681) );
  INV_X1 U3960 ( .A(n1003), .ZN(n3682) );
  NOR2_X1 U3961 ( .A1(n1431), .A2(n1458), .ZN(n777) );
  NAND2_X1 U3962 ( .A1(n3703), .A2(n778), .ZN(n558) );
  OAI22_X1 U3963 ( .A1(n434), .A2(n3005), .B1(n3004), .B2(n384), .ZN(n2442) );
  BUF_X1 U3964 ( .A(n3553), .Z(n3684) );
  BUF_X1 U3965 ( .A(n781), .Z(n3685) );
  INV_X1 U3966 ( .A(n3468), .ZN(n876) );
  OAI21_X1 U3967 ( .B1(n3568), .B2(n3741), .A(n3438), .ZN(n2434) );
  AOI21_X2 U3968 ( .B1(n878), .B2(n897), .A(n879), .ZN(n877) );
  AOI21_X2 U3969 ( .B1(n885), .B2(n893), .A(n886), .ZN(n884) );
  OAI21_X1 U3970 ( .B1(n884), .B2(n880), .A(n881), .ZN(n879) );
  INV_X1 U3971 ( .A(n814), .ZN(n1011) );
  OAI21_X1 U3972 ( .B1(n816), .B2(n814), .A(n815), .ZN(n813) );
  NOR2_X2 U3973 ( .A1(n1642), .A2(n1669), .ZN(n814) );
  OAI22_X1 U3974 ( .A1(n437), .A2(n2979), .B1(n2978), .B2(n387), .ZN(n2415) );
  NAND2_X1 U3975 ( .A1(n809), .A2(n817), .ZN(n807) );
  INV_X1 U3976 ( .A(n706), .ZN(n3688) );
  INV_X1 U3977 ( .A(n3688), .ZN(n3689) );
  OAI22_X1 U3978 ( .A1(n434), .A2(n3012), .B1(n3011), .B2(n384), .ZN(n2449) );
  OAI21_X1 U3979 ( .B1(n896), .B2(n883), .A(n884), .ZN(n882) );
  NAND2_X2 U3980 ( .A1(n1918), .A2(n1933), .ZN(n888) );
  NAND2_X2 U3981 ( .A1(n1519), .A2(n1550), .ZN(n794) );
  XOR2_X2 U3982 ( .A(n3472), .B(a[6]), .Z(n3691) );
  XNOR2_X1 U3983 ( .A(n749), .B(n553), .ZN(product[42]) );
  INV_X1 U3984 ( .A(n793), .ZN(n791) );
  AOI21_X1 U3985 ( .B1(n795), .B2(n791), .A(n792), .ZN(n790) );
  XNOR2_X1 U3986 ( .A(n795), .B(n561), .ZN(product[34]) );
  NAND2_X1 U3987 ( .A1(n1553), .A2(n1583), .ZN(n3692) );
  NAND2_X1 U3988 ( .A1(n1553), .A2(n1555), .ZN(n3693) );
  NAND2_X1 U3989 ( .A1(n1583), .A2(n1555), .ZN(n3694) );
  NAND3_X1 U3990 ( .A1(n3692), .A2(n3694), .A3(n3693), .ZN(n1550) );
  NOR2_X1 U3991 ( .A1(n428), .A2(n3077), .ZN(n3696) );
  NOR2_X1 U3992 ( .A1(n3076), .A2(n3639), .ZN(n3697) );
  XNOR2_X1 U3993 ( .A(n503), .B(n330), .ZN(n3077) );
  INV_X1 U3994 ( .A(n3560), .ZN(n1003) );
  OR2_X1 U3995 ( .A1(n1377), .A2(n1402), .ZN(n3698) );
  OAI21_X1 U3996 ( .B1(n3672), .B2(n3691), .A(n330), .ZN(n2502) );
  OAI21_X1 U3997 ( .B1(n800), .B2(n804), .A(n801), .ZN(n3699) );
  BUF_X1 U3998 ( .A(n612), .Z(n3700) );
  INV_X1 U3999 ( .A(n3579), .ZN(n855) );
  NAND2_X1 U4000 ( .A1(n3480), .A2(n3456), .ZN(n569) );
  NOR2_X1 U4001 ( .A1(n446), .A2(n2885), .ZN(n3701) );
  NOR2_X1 U4002 ( .A1(n2884), .A2(n396), .ZN(n3702) );
  OR2_X1 U4003 ( .A1(n3701), .A2(n3702), .ZN(n2318) );
  XNOR2_X1 U4004 ( .A(n491), .B(n348), .ZN(n2885) );
  XOR2_X1 U4005 ( .A(n3695), .B(n348), .Z(n3234) );
  NAND2_X1 U4006 ( .A1(n1670), .A2(n1697), .ZN(n820) );
  NAND2_X1 U4007 ( .A1(n1377), .A2(n1402), .ZN(n770) );
  NAND2_X1 U4008 ( .A1(n786), .A2(n798), .ZN(n784) );
  OR2_X1 U4009 ( .A1(n3681), .A2(n1458), .ZN(n3703) );
  XNOR2_X1 U4010 ( .A(n1520), .B(n1493), .ZN(n3704) );
  BUF_X1 U4011 ( .A(n3528), .Z(n3705) );
  INV_X1 U4012 ( .A(n861), .ZN(n1018) );
  NAND2_X1 U4013 ( .A1(n775), .A2(n3512), .ZN(n765) );
  INV_X1 U4014 ( .A(n794), .ZN(n792) );
  NAND2_X1 U4015 ( .A1(n791), .A2(n794), .ZN(n561) );
  NOR2_X1 U4016 ( .A1(n3684), .A2(n1488), .ZN(n3706) );
  NOR2_X1 U4017 ( .A1(n3542), .A2(n3068), .ZN(n3707) );
  NOR2_X1 U4018 ( .A1(n3067), .A2(n3639), .ZN(n3708) );
  XNOR2_X1 U4019 ( .A(n521), .B(n330), .ZN(n3068) );
  XNOR2_X1 U4020 ( .A(n523), .B(n330), .ZN(n3067) );
  NAND2_X1 U4021 ( .A1(n1820), .A2(n1841), .ZN(n862) );
  NOR2_X1 U4022 ( .A1(n446), .A2(n2884), .ZN(n3710) );
  NOR2_X1 U4023 ( .A1(n2883), .A2(n396), .ZN(n3711) );
  OR2_X1 U4024 ( .A1(n3710), .A2(n3711), .ZN(n2317) );
  XNOR2_X1 U4025 ( .A(n493), .B(n348), .ZN(n2884) );
  NOR2_X2 U4026 ( .A1(n1519), .A2(n1550), .ZN(n793) );
  NOR2_X1 U4027 ( .A1(n452), .A2(n2818), .ZN(n3713) );
  NOR2_X1 U4028 ( .A1(n2817), .A2(n402), .ZN(n3714) );
  XNOR2_X1 U4029 ( .A(n493), .B(n354), .ZN(n2818) );
  XNOR2_X1 U4030 ( .A(n495), .B(n354), .ZN(n2817) );
  NAND2_X1 U4031 ( .A1(n1759), .A2(n1736), .ZN(n3715) );
  NAND2_X1 U4032 ( .A1(n1759), .A2(n1738), .ZN(n3716) );
  NAND2_X1 U4033 ( .A1(n1736), .A2(n1738), .ZN(n3717) );
  NAND3_X1 U4034 ( .A1(n3715), .A2(n3717), .A3(n3716), .ZN(n1729) );
  XOR2_X1 U4035 ( .A(n3718), .B(n330), .Z(n3240) );
  NAND2_X1 U4036 ( .A1(n686), .A2(n673), .ZN(n671) );
  NAND2_X1 U4037 ( .A1(n1005), .A2(n781), .ZN(n559) );
  OAI21_X1 U4038 ( .B1(n728), .B2(n613), .A(n614), .ZN(n612) );
  NAND2_X1 U4039 ( .A1(n1491), .A2(n1520), .ZN(n3719) );
  NAND2_X1 U4040 ( .A1(n1491), .A2(n1493), .ZN(n3720) );
  NAND2_X1 U4041 ( .A1(n1520), .A2(n1493), .ZN(n3721) );
  NAND3_X1 U4042 ( .A1(n3719), .A2(n3721), .A3(n3720), .ZN(n1488) );
  NOR2_X1 U4043 ( .A1(n446), .A2(n2883), .ZN(n3722) );
  NOR2_X1 U4044 ( .A1(n2882), .A2(n396), .ZN(n3723) );
  OR2_X1 U4045 ( .A1(n3722), .A2(n3723), .ZN(n2316) );
  XNOR2_X1 U4046 ( .A(n495), .B(n348), .ZN(n2883) );
  XNOR2_X1 U4047 ( .A(n497), .B(n348), .ZN(n2882) );
  AND2_X2 U4048 ( .A1(n3237), .A2(n3540), .ZN(n3724) );
  BUF_X8 U4049 ( .A(n3479), .Z(n3726) );
  INV_X1 U4050 ( .A(n3481), .ZN(n1010) );
  NAND2_X1 U4051 ( .A1(n1612), .A2(n1641), .ZN(n812) );
  OAI22_X1 U4052 ( .A1(n3435), .A2(n2983), .B1(n2982), .B2(n387), .ZN(n2419)
         );
  NAND2_X1 U4053 ( .A1(n844), .A2(n847), .ZN(n570) );
  NAND2_X2 U4054 ( .A1(n844), .A2(n851), .ZN(n842) );
  NOR2_X2 U4055 ( .A1(n1774), .A2(n1797), .ZN(n846) );
  NAND2_X1 U4056 ( .A1(n1774), .A2(n1797), .ZN(n847) );
  NAND2_X1 U4057 ( .A1(n1750), .A2(n1773), .ZN(n840) );
  NOR2_X2 U4058 ( .A1(n765), .A2(n784), .ZN(n763) );
  INV_X1 U4059 ( .A(n3602), .ZN(n3759) );
  OAI21_X1 U4060 ( .B1(n3669), .B2(n773), .A(n770), .ZN(n768) );
  BUF_X1 U4061 ( .A(n603), .Z(n3732) );
  NOR2_X1 U4062 ( .A1(n446), .A2(n2880), .ZN(n3733) );
  NOR2_X1 U4063 ( .A1(n2879), .A2(n396), .ZN(n3734) );
  XNOR2_X1 U4064 ( .A(n501), .B(n348), .ZN(n2880) );
  XNOR2_X1 U4065 ( .A(n503), .B(n348), .ZN(n2879) );
  NAND2_X1 U4066 ( .A1(n832), .A2(n838), .ZN(n3735) );
  INV_X1 U4067 ( .A(n833), .ZN(n3736) );
  NOR2_X1 U4068 ( .A1(n3542), .A2(n3076), .ZN(n3737) );
  NOR2_X1 U4069 ( .A1(n3075), .A2(n3639), .ZN(n3738) );
  INV_X2 U4070 ( .A(n3739), .ZN(n3740) );
  NOR2_X2 U4071 ( .A1(n830), .A2(n842), .ZN(n828) );
  INV_X1 U4072 ( .A(n835), .ZN(n833) );
  XNOR2_X1 U4073 ( .A(n505), .B(n330), .ZN(n3076) );
  XNOR2_X1 U4074 ( .A(n507), .B(n330), .ZN(n3075) );
  AND2_X2 U4075 ( .A1(n3238), .A2(n384), .ZN(n3741) );
  INV_X4 U4076 ( .A(n3741), .ZN(n434) );
  INV_X1 U4077 ( .A(n3490), .ZN(n797) );
  NAND2_X2 U4078 ( .A1(n1582), .A2(n1611), .ZN(n804) );
  NAND2_X2 U4079 ( .A1(n1281), .A2(n1302), .ZN(n739) );
  NAND2_X1 U4080 ( .A1(n832), .A2(n835), .ZN(n568) );
  INV_X1 U4081 ( .A(n3650), .ZN(n3758) );
  XNOR2_X1 U4082 ( .A(n650), .B(n539), .ZN(product[56]) );
  XNOR2_X1 U4083 ( .A(n643), .B(n538), .ZN(product[57]) );
  INV_X1 U4084 ( .A(n3727), .ZN(n826) );
  XNOR2_X1 U4085 ( .A(n737), .B(n551), .ZN(product[44]) );
  XOR2_X1 U4086 ( .A(n665), .B(n542), .Z(product[53]) );
  AOI21_X2 U4087 ( .B1(n3621), .B2(n989), .A(n667), .ZN(n665) );
  INV_X1 U4088 ( .A(n783), .ZN(n782) );
  OAI21_X1 U4089 ( .B1(n774), .B2(n3682), .A(n3585), .ZN(n771) );
  XOR2_X1 U4090 ( .A(n774), .B(n557), .Z(product[38]) );
  OAI21_X2 U4091 ( .B1(n630), .B2(n624), .A(n625), .ZN(n623) );
  XOR2_X1 U4092 ( .A(n630), .B(n537), .Z(product[58]) );
  INV_X1 U4093 ( .A(n683), .ZN(n682) );
  AOI21_X2 U4094 ( .B1(n683), .B2(n631), .A(n632), .ZN(n630) );
  OAI21_X1 U4095 ( .B1(n744), .B2(n738), .A(n739), .ZN(n737) );
  INV_X1 U4096 ( .A(n3505), .ZN(n1006) );
  XNOR2_X1 U4097 ( .A(n3689), .B(n548), .ZN(product[47]) );
  AOI21_X2 U4098 ( .B1(n706), .B2(n994), .A(n703), .ZN(n701) );
  XNOR2_X1 U4099 ( .A(n761), .B(n555), .ZN(product[40]) );
  OAI21_X1 U4100 ( .B1(n724), .B2(n718), .A(n719), .ZN(n717) );
  XOR2_X1 U4101 ( .A(n724), .B(n550), .Z(product[45]) );
  AOI21_X1 U4102 ( .B1(n761), .B2(n757), .A(n758), .ZN(n756) );
  AOI21_X1 U4103 ( .B1(n761), .B2(n611), .A(n3700), .ZN(n610) );
  AOI21_X2 U4104 ( .B1(n761), .B2(n3485), .A(n726), .ZN(n724) );
  XOR2_X1 U4105 ( .A(n3551), .B(n552), .Z(product[43]) );
  NAND2_X1 U4106 ( .A1(n3681), .A2(n1458), .ZN(n778) );
  OAI21_X1 U4107 ( .B1(n782), .B2(n3706), .A(n3685), .ZN(n779) );
  INV_X1 U4108 ( .A(n3706), .ZN(n1005) );
  INV_X1 U4109 ( .A(n3538), .ZN(n3756) );
  XOR2_X1 U4110 ( .A(n3648), .B(n533), .Z(product[62]) );
  OAI21_X1 U4111 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  INV_X8 U4112 ( .A(n3751), .ZN(n381) );
  XNOR2_X1 U4113 ( .A(n670), .B(n543), .ZN(product[52]) );
  OAI21_X1 U4114 ( .B1(n3545), .B2(n651), .A(n652), .ZN(n650) );
  OAI21_X1 U4115 ( .B1(n653), .B2(n644), .A(n645), .ZN(n643) );
  XOR2_X1 U4116 ( .A(n3546), .B(n540), .Z(product[55]) );
  XNOR2_X1 U4117 ( .A(n3732), .B(n534), .ZN(product[61]) );
  INV_X1 U4118 ( .A(n3670), .ZN(n761) );
  INV_X2 U4119 ( .A(n594), .ZN(product[1]) );
  INV_X2 U4120 ( .A(n699), .ZN(n993) );
  INV_X2 U4121 ( .A(n696), .ZN(n992) );
  INV_X2 U4122 ( .A(n680), .ZN(n991) );
  INV_X2 U4123 ( .A(n677), .ZN(n990) );
  INV_X2 U4124 ( .A(n663), .ZN(n988) );
  INV_X2 U4125 ( .A(n660), .ZN(n987) );
  INV_X2 U4126 ( .A(n651), .ZN(n986) );
  INV_X2 U4127 ( .A(n648), .ZN(n985) );
  INV_X2 U4128 ( .A(n596), .ZN(n979) );
  INV_X2 U4129 ( .A(n978), .ZN(n976) );
  INV_X2 U4130 ( .A(n975), .ZN(n973) );
  INV_X2 U4131 ( .A(n967), .ZN(n965) );
  INV_X2 U4132 ( .A(n959), .ZN(n957) );
  INV_X2 U4133 ( .A(n955), .ZN(n954) );
  INV_X2 U4134 ( .A(n953), .ZN(n951) );
  INV_X2 U4135 ( .A(n948), .ZN(n946) );
  INV_X2 U4136 ( .A(n941), .ZN(n939) );
  INV_X2 U4137 ( .A(n937), .ZN(n936) );
  INV_X2 U4138 ( .A(n935), .ZN(n933) );
  INV_X2 U4139 ( .A(n930), .ZN(n928) );
  INV_X2 U4140 ( .A(n924), .ZN(n923) );
  INV_X2 U4141 ( .A(n915), .ZN(n914) );
  INV_X2 U4142 ( .A(n913), .ZN(n911) );
  INV_X2 U4143 ( .A(n903), .ZN(n901) );
  INV_X2 U4144 ( .A(n897), .ZN(n896) );
  INV_X2 U4145 ( .A(n891), .ZN(n893) );
  INV_X2 U4146 ( .A(n888), .ZN(n886) );
  INV_X2 U4147 ( .A(n875), .ZN(n873) );
  INV_X2 U4148 ( .A(n840), .ZN(n838) );
  INV_X2 U4149 ( .A(n748), .ZN(n746) );
  INV_X2 U4150 ( .A(n747), .ZN(n999) );
  INV_X2 U4151 ( .A(n736), .ZN(n734) );
  INV_X2 U4152 ( .A(n735), .ZN(n997) );
  INV_X2 U4153 ( .A(n719), .ZN(n721) );
  INV_X2 U4154 ( .A(n718), .ZN(n996) );
  INV_X2 U4155 ( .A(n716), .ZN(n714) );
  INV_X2 U4156 ( .A(n715), .ZN(n995) );
  INV_X2 U4157 ( .A(n712), .ZN(n710) );
  INV_X2 U4158 ( .A(n711), .ZN(n709) );
  INV_X2 U4159 ( .A(n705), .ZN(n703) );
  INV_X2 U4160 ( .A(n704), .ZN(n994) );
  INV_X2 U4161 ( .A(n691), .ZN(n689) );
  INV_X2 U4162 ( .A(n690), .ZN(n688) );
  INV_X2 U4163 ( .A(n669), .ZN(n667) );
  INV_X2 U4164 ( .A(n668), .ZN(n989) );
  INV_X2 U4165 ( .A(n657), .ZN(n655) );
  INV_X2 U4166 ( .A(n656), .ZN(n654) );
  INV_X2 U4167 ( .A(n647), .ZN(n645) );
  INV_X2 U4168 ( .A(n646), .ZN(n644) );
  INV_X2 U4169 ( .A(n642), .ZN(n640) );
  INV_X2 U4170 ( .A(n641), .ZN(n984) );
  INV_X2 U4171 ( .A(n633), .ZN(n631) );
  INV_X2 U4172 ( .A(n625), .ZN(n627) );
  INV_X2 U4173 ( .A(n624), .ZN(n983) );
  INV_X2 U4174 ( .A(n622), .ZN(n620) );
  INV_X2 U4175 ( .A(n621), .ZN(n982) );
  INV_X2 U4176 ( .A(n609), .ZN(n607) );
  INV_X2 U4177 ( .A(n608), .ZN(n981) );
  INV_X2 U4178 ( .A(n602), .ZN(n600) );
  INV_X2 U4179 ( .A(n601), .ZN(n980) );
  INV_X2 U4180 ( .A(n3578), .ZN(n3292) );
  INV_X2 U4181 ( .A(n3726), .ZN(n3290) );
  INV_X2 U4182 ( .A(n3531), .ZN(n3288) );
  INV_X2 U4183 ( .A(n3438), .ZN(n3287) );
  INV_X2 U4184 ( .A(n3712), .ZN(n3284) );
  INV_X2 U4185 ( .A(n348), .ZN(n3283) );
  INV_X2 U4186 ( .A(n357), .ZN(n3280) );
  INV_X2 U4187 ( .A(n360), .ZN(n3279) );
  INV_X2 U4188 ( .A(n363), .ZN(n3278) );
  NAND2_X2 U4189 ( .A1(n3578), .A2(n3440), .ZN(n3195) );
  NAND2_X2 U4190 ( .A1(n324), .A2(n3440), .ZN(n3162) );
  NAND2_X2 U4191 ( .A1(n3740), .A2(n3440), .ZN(n3129) );
  NAND2_X2 U4192 ( .A1(n330), .A2(n3440), .ZN(n3096) );
  NAND2_X2 U4193 ( .A1(n3531), .A2(n3440), .ZN(n3063) );
  NAND2_X2 U4194 ( .A1(n3438), .A2(n3440), .ZN(n3030) );
  NAND2_X2 U4195 ( .A1(n339), .A2(n3440), .ZN(n2997) );
  NAND2_X2 U4196 ( .A1(n342), .A2(n3440), .ZN(n2964) );
  NAND2_X2 U4197 ( .A1(n3712), .A2(n3440), .ZN(n2931) );
  NAND2_X2 U4198 ( .A1(n348), .A2(n3440), .ZN(n2898) );
  NAND2_X2 U4199 ( .A1(n351), .A2(n3440), .ZN(n2865) );
  NAND2_X2 U4200 ( .A1(n3605), .A2(n3440), .ZN(n2832) );
  NAND2_X2 U4201 ( .A1(n357), .A2(n3440), .ZN(n2799) );
  NAND2_X2 U4202 ( .A1(n360), .A2(n3440), .ZN(n2766) );
  NAND2_X2 U4203 ( .A1(n363), .A2(n3440), .ZN(n2733) );
  NAND2_X2 U4204 ( .A1(n366), .A2(n3440), .ZN(n2700) );
  NOR2_X2 U4205 ( .A1(n3425), .A2(n3440), .ZN(n2603) );
  NOR2_X2 U4206 ( .A1(n375), .A2(n3440), .ZN(n2569) );
  NOR2_X2 U4207 ( .A1(n381), .A2(n3440), .ZN(n2501) );
  NOR2_X2 U4208 ( .A1(n384), .A2(n3440), .ZN(n2467) );
  NOR2_X2 U4209 ( .A1(n387), .A2(n3440), .ZN(n2433) );
  NOR2_X2 U4210 ( .A1(n390), .A2(n3440), .ZN(n2399) );
  NOR2_X2 U4211 ( .A1(n3556), .A2(n3440), .ZN(n2365) );
  NOR2_X2 U4212 ( .A1(n396), .A2(n3440), .ZN(n2331) );
  NOR2_X2 U4213 ( .A1(n399), .A2(n3440), .ZN(n2297) );
  NOR2_X2 U4214 ( .A1(n402), .A2(n3440), .ZN(n2263) );
  NOR2_X2 U4215 ( .A1(n3460), .A2(n3440), .ZN(n2229) );
  NOR2_X2 U4216 ( .A1(n408), .A2(n3440), .ZN(n2195) );
  NOR2_X2 U4217 ( .A1(n3557), .A2(n3440), .ZN(n2161) );
  INV_X2 U4218 ( .A(n1548), .ZN(n1580) );
  INV_X2 U4219 ( .A(n1486), .ZN(n1487) );
  INV_X2 U4220 ( .A(n1374), .ZN(n1375) );
  INV_X2 U4221 ( .A(n1324), .ZN(n1325) );
  INV_X2 U4222 ( .A(n1278), .ZN(n1279) );
  INV_X2 U4223 ( .A(n1236), .ZN(n1237) );
  INV_X2 U4224 ( .A(n1198), .ZN(n1199) );
  INV_X2 U4225 ( .A(n1164), .ZN(n1165) );
  INV_X2 U4226 ( .A(n1134), .ZN(n1135) );
  INV_X2 U4227 ( .A(n1108), .ZN(n1109) );
  INV_X2 U4228 ( .A(n1086), .ZN(n1087) );
  INV_X2 U4229 ( .A(n1068), .ZN(n1069) );
  INV_X2 U4230 ( .A(n1054), .ZN(n1055) );
  INV_X2 U4231 ( .A(n1044), .ZN(n1045) );
  XOR2_X1 U4232 ( .A(n3760), .B(n3761), .Z(n1041) );
  XOR2_X1 U4233 ( .A(n2077), .B(n1044), .Z(n3761) );
  INV_X2 U4234 ( .A(n977), .ZN(n1040) );
  INV_X2 U4235 ( .A(n974), .ZN(n972) );
  INV_X2 U4236 ( .A(n969), .ZN(n1038) );
  INV_X2 U4237 ( .A(n966), .ZN(n964) );
  INV_X2 U4238 ( .A(n961), .ZN(n1036) );
  INV_X2 U4239 ( .A(n958), .ZN(n956) );
  INV_X2 U4240 ( .A(n952), .ZN(n950) );
  INV_X2 U4241 ( .A(n947), .ZN(n945) );
  INV_X2 U4242 ( .A(n940), .ZN(n938) );
  INV_X2 U4243 ( .A(n934), .ZN(n932) );
  INV_X2 U4244 ( .A(n929), .ZN(n927) );
  INV_X2 U4245 ( .A(n921), .ZN(n1029) );
  INV_X2 U4246 ( .A(n918), .ZN(n1028) );
  INV_X2 U4247 ( .A(n912), .ZN(n910) );
  INV_X2 U4248 ( .A(n902), .ZN(n900) );
  INV_X2 U4249 ( .A(n890), .ZN(n892) );
  INV_X2 U4250 ( .A(n887), .ZN(n885) );
  INV_X2 U4251 ( .A(n880), .ZN(n1022) );
  INV_X2 U4252 ( .A(n874), .ZN(n872) );
  INV_X2 U4253 ( .A(n869), .ZN(n1020) );
  INV_X2 U4254 ( .A(n864), .ZN(n1019) );
  INV_X2 U4255 ( .A(n849), .ZN(n851) );
  INV_X2 U4256 ( .A(n846), .ZN(n844) );
  INV_X2 U4257 ( .A(n824), .ZN(n822) );
  INV_X2 U4258 ( .A(n759), .ZN(n757) );
endmodule


module reg64_2 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  DFFR_X2 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X2 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X2 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module reg64_1 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  DFFR_X1 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  DFFR_X2 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  DFFR_X2 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X2 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X2 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module reg64_0 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  DFFR_X2 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X2 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X1 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module mul32_2 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_2_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module mul32_1 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_1_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module mul32_0 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_0_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module reg64_3 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  DFFR_X1 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  DFFR_X1 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X2 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module mul32_3 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_3_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module mulcascade ( a0, b0, a1, b1, a2, b2, a3, b3, result0, result1, result2, 
        result3, resetn, clk );
  input [31:0] a0;
  input [31:0] b0;
  input [31:0] a1;
  input [31:0] b1;
  input [31:0] a2;
  input [31:0] b2;
  input [31:0] a3;
  input [31:0] b3;
  output [63:0] result0;
  output [63:0] result1;
  output [63:0] result2;
  output [63:0] result3;
  input resetn, clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269;
  wire   [63:0] reg0in;
  wire   [63:0] reg1in;
  wire   [63:0] reg2in;
  wire   [63:0] reg3in;

  mul32_3 mul0 ( .a({a0[31], n8, a0[29], n18, a0[27:23], n14, a0[21], n4, 
        a0[19:11], n2, a0[9], n10, a0[7:0]}), .b({n158, n170, n180, n164, n168, 
        n174, n152, n154, n196, n142, n266, n264, n254, n260, n250, n238, n248, 
        n244, n234, n222, n232, n228, n218, n206, n216, n212, n202, n190, n200, 
        n186, n184, b0[0]}), .result(reg0in) );
  reg64_3 reg0 ( .d(reg0in), .resetn(n269), .clk(clk), .q(result0) );
  mul32_2 mul1 ( .a({a1[31:17], n6, a1[15:3], n16, a1[1:0]}), .b({n148, n138, 
        n136, n132, n126, n122, n116, n120, n110, n106, n100, n104, n94, n90, 
        n84, n88, n78, n74, n68, n72, n62, n58, n52, n56, n46, n42, n36, n40, 
        n30, n26, n24, b1[0]}), .result(reg1in) );
  reg64_2 reg1 ( .d(reg1in), .resetn(n269), .clk(clk), .q(result1) );
  mul32_1 mul2 ( .a({a2[31:19], n12, a2[17], n20, a2[15:0]}), .b({n50, n60, 
        n70, n76, n82, n86, n96, n92, n98, n102, n112, n108, n114, n118, n128, 
        n124, n130, n134, n144, n140, n146, n150, n160, n156, n162, n166, n176, 
        n172, n178, n182, n192, b2[0]}), .result(reg2in) );
  reg64_1 reg2 ( .d(reg2in), .resetn(n269), .clk(clk), .q(result2) );
  mul32_0 mul3 ( .a(a3), .b({n204, n214, n226, n230, n242, n246, n252, n262, 
        n32, n22, n268, n38, n28, n258, n44, n34, n256, n54, n48, n240, n64, 
        n188, n236, n66, n194, n224, n80, n198, n220, n210, n208, b3[0]}), 
        .result(reg3in) );
  reg64_0 reg4 ( .d(reg3in), .resetn(n269), .clk(clk), .q(result3) );
  INV_X1 U1 ( .A(b2[2]), .ZN(n181) );
  INV_X1 U2 ( .A(a0[28]), .ZN(n17) );
  INV_X1 U3 ( .A(a0[20]), .ZN(n3) );
  INV_X1 U4 ( .A(b2[10]), .ZN(n149) );
  INV_X1 U5 ( .A(b2[6]), .ZN(n165) );
  INV_X1 U6 ( .A(a0[30]), .ZN(n7) );
  INV_X1 U7 ( .A(b1[11]), .ZN(n61) );
  INV_X1 U8 ( .A(b2[18]), .ZN(n117) );
  INV_X1 U9 ( .A(b2[14]), .ZN(n133) );
  INV_X1 U10 ( .A(a0[8]), .ZN(n9) );
  INV_X1 U11 ( .A(a1[16]), .ZN(n5) );
  INV_X1 U12 ( .A(b2[22]), .ZN(n101) );
  INV_X1 U13 ( .A(a0[22]), .ZN(n13) );
  INV_X1 U14 ( .A(a2[18]), .ZN(n11) );
  INV_X1 U15 ( .A(b1[2]), .ZN(n25) );
  INV_X1 U16 ( .A(b3[22]), .ZN(n21) );
  INV_X1 U17 ( .A(b2[29]), .ZN(n69) );
  INV_X1 U18 ( .A(b2[26]), .ZN(n85) );
  INV_X1 U19 ( .A(b1[5]), .ZN(n35) );
  INV_X1 U20 ( .A(b1[7]), .ZN(n45) );
  INV_X1 U21 ( .A(b3[14]), .ZN(n53) );
  INV_X1 U22 ( .A(b1[3]), .ZN(n29) );
  INV_X1 U23 ( .A(b3[16]), .ZN(n33) );
  INV_X1 U24 ( .A(b3[20]), .ZN(n37) );
  INV_X1 U25 ( .A(b3[23]), .ZN(n31) );
  INV_X1 U26 ( .A(b1[1]), .ZN(n23) );
  INV_X1 U27 ( .A(b1[6]), .ZN(n41) );
  INV_X1 U28 ( .A(b3[19]), .ZN(n27) );
  INV_X1 U29 ( .A(b2[31]), .ZN(n49) );
  INV_X1 U30 ( .A(b1[4]), .ZN(n39) );
  INV_X1 U31 ( .A(b3[17]), .ZN(n43) );
  INV_X1 U32 ( .A(b3[13]), .ZN(n47) );
  INV_X1 U33 ( .A(b1[9]), .ZN(n51) );
  INV_X1 U34 ( .A(b2[30]), .ZN(n59) );
  INV_X1 U35 ( .A(b1[10]), .ZN(n57) );
  INV_X1 U36 ( .A(b1[13]), .ZN(n67) );
  INV_X1 U37 ( .A(b3[8]), .ZN(n65) );
  INV_X1 U38 ( .A(b1[14]), .ZN(n73) );
  INV_X1 U39 ( .A(b1[8]), .ZN(n55) );
  INV_X1 U40 ( .A(b3[11]), .ZN(n63) );
  INV_X1 U41 ( .A(b1[12]), .ZN(n71) );
  INV_X1 U42 ( .A(b2[28]), .ZN(n75) );
  INV_X1 U43 ( .A(b1[17]), .ZN(n83) );
  INV_X1 U44 ( .A(b2[27]), .ZN(n81) );
  INV_X1 U45 ( .A(b2[24]), .ZN(n91) );
  INV_X1 U46 ( .A(b1[18]), .ZN(n89) );
  INV_X1 U47 ( .A(b3[5]), .ZN(n79) );
  INV_X1 U48 ( .A(b1[22]), .ZN(n105) );
  INV_X1 U49 ( .A(b1[16]), .ZN(n87) );
  INV_X1 U50 ( .A(b1[21]), .ZN(n99) );
  INV_X1 U51 ( .A(b2[23]), .ZN(n97) );
  INV_X1 U52 ( .A(b1[20]), .ZN(n103) );
  INV_X1 U53 ( .A(b2[20]), .ZN(n107) );
  INV_X1 U54 ( .A(b2[19]), .ZN(n113) );
  INV_X1 U55 ( .A(b2[25]), .ZN(n95) );
  INV_X1 U56 ( .A(b2[16]), .ZN(n123) );
  INV_X1 U57 ( .A(b1[26]), .ZN(n121) );
  INV_X1 U58 ( .A(b2[21]), .ZN(n111) );
  INV_X1 U59 ( .A(b1[25]), .ZN(n115) );
  INV_X1 U60 ( .A(b1[30]), .ZN(n137) );
  INV_X1 U61 ( .A(b1[24]), .ZN(n119) );
  INV_X1 U62 ( .A(b1[28]), .ZN(n131) );
  INV_X1 U63 ( .A(b2[15]), .ZN(n129) );
  INV_X1 U64 ( .A(b1[29]), .ZN(n135) );
  INV_X1 U65 ( .A(b2[12]), .ZN(n139) );
  INV_X1 U66 ( .A(b2[11]), .ZN(n145) );
  INV_X1 U67 ( .A(b2[17]), .ZN(n127) );
  INV_X1 U68 ( .A(b2[8]), .ZN(n155) );
  INV_X1 U69 ( .A(b0[24]), .ZN(n153) );
  INV_X1 U70 ( .A(b2[13]), .ZN(n143) );
  INV_X1 U71 ( .A(b1[31]), .ZN(n147) );
  INV_X1 U72 ( .A(b0[30]), .ZN(n169) );
  INV_X1 U73 ( .A(b0[25]), .ZN(n151) );
  INV_X1 U74 ( .A(b0[28]), .ZN(n163) );
  INV_X1 U75 ( .A(b2[7]), .ZN(n161) );
  INV_X1 U76 ( .A(b2[4]), .ZN(n171) );
  INV_X1 U77 ( .A(b2[3]), .ZN(n177) );
  INV_X1 U78 ( .A(b2[9]), .ZN(n159) );
  INV_X1 U79 ( .A(b0[2]), .ZN(n185) );
  INV_X1 U80 ( .A(b0[27]), .ZN(n167) );
  INV_X1 U81 ( .A(b2[5]), .ZN(n175) );
  INV_X1 U82 ( .A(b0[29]), .ZN(n179) );
  INV_X1 U83 ( .A(b3[10]), .ZN(n187) );
  INV_X1 U84 ( .A(b0[23]), .ZN(n195) );
  INV_X1 U85 ( .A(b3[7]), .ZN(n193) );
  INV_X1 U86 ( .A(b0[5]), .ZN(n201) );
  INV_X1 U87 ( .A(b0[1]), .ZN(n183) );
  INV_X1 U88 ( .A(b3[2]), .ZN(n209) );
  INV_X1 U89 ( .A(b2[1]), .ZN(n191) );
  INV_X1 U90 ( .A(b0[3]), .ZN(n199) );
  INV_X1 U91 ( .A(b3[31]), .ZN(n203) );
  INV_X1 U92 ( .A(b3[1]), .ZN(n207) );
  INV_X1 U93 ( .A(b0[6]), .ZN(n211) );
  INV_X1 U94 ( .A(b3[3]), .ZN(n219) );
  INV_X1 U95 ( .A(b0[9]), .ZN(n217) );
  INV_X1 U96 ( .A(b0[10]), .ZN(n227) );
  INV_X1 U97 ( .A(b3[29]), .ZN(n225) );
  INV_X1 U98 ( .A(b0[7]), .ZN(n215) );
  INV_X1 U99 ( .A(b3[27]), .ZN(n241) );
  INV_X1 U100 ( .A(b3[6]), .ZN(n223) );
  INV_X1 U101 ( .A(b3[9]), .ZN(n235) );
  INV_X1 U102 ( .A(b0[13]), .ZN(n233) );
  INV_X1 U103 ( .A(b3[12]), .ZN(n239) );
  INV_X1 U104 ( .A(b0[14]), .ZN(n243) );
  INV_X1 U105 ( .A(b0[11]), .ZN(n231) );
  INV_X1 U106 ( .A(b0[18]), .ZN(n259) );
  INV_X1 U107 ( .A(b3[18]), .ZN(n257) );
  INV_X1 U108 ( .A(b3[25]), .ZN(n251) );
  INV_X1 U109 ( .A(b0[17]), .ZN(n249) );
  INV_X1 U110 ( .A(b3[15]), .ZN(n255) );
  INV_X1 U111 ( .A(b0[15]), .ZN(n247) );
  INV_X1 U112 ( .A(b0[16]), .ZN(n237) );
  INV_X1 U113 ( .A(b0[19]), .ZN(n253) );
  INV_X1 U114 ( .A(b0[21]), .ZN(n265) );
  INV_X1 U115 ( .A(b0[8]), .ZN(n205) );
  INV_X1 U116 ( .A(b0[12]), .ZN(n221) );
  INV_X1 U117 ( .A(b0[20]), .ZN(n263) );
  INV_X1 U118 ( .A(b3[21]), .ZN(n267) );
  INV_X1 U119 ( .A(b0[26]), .ZN(n173) );
  INV_X1 U120 ( .A(b0[4]), .ZN(n189) );
  INV_X1 U121 ( .A(b3[24]), .ZN(n261) );
  BUF_X1 U122 ( .A(resetn), .Z(n269) );
  INV_X1 U123 ( .A(b0[22]), .ZN(n141) );
  INV_X1 U124 ( .A(b0[31]), .ZN(n157) );
  INV_X1 U125 ( .A(b3[28]), .ZN(n229) );
  INV_X1 U126 ( .A(b3[26]), .ZN(n245) );
  INV_X1 U127 ( .A(b1[23]), .ZN(n109) );
  INV_X1 U128 ( .A(b1[27]), .ZN(n125) );
  INV_X1 U129 ( .A(b3[4]), .ZN(n197) );
  INV_X1 U130 ( .A(b3[30]), .ZN(n213) );
  INV_X1 U131 ( .A(b1[15]), .ZN(n77) );
  INV_X1 U132 ( .A(b1[19]), .ZN(n93) );
  INV_X1 U133 ( .A(a0[10]), .ZN(n1) );
  INV_X1 U134 ( .A(n1), .ZN(n2) );
  INV_X1 U135 ( .A(n3), .ZN(n4) );
  INV_X1 U136 ( .A(n5), .ZN(n6) );
  INV_X1 U137 ( .A(n7), .ZN(n8) );
  INV_X1 U138 ( .A(n9), .ZN(n10) );
  INV_X1 U139 ( .A(n11), .ZN(n12) );
  INV_X1 U140 ( .A(n13), .ZN(n14) );
  INV_X4 U141 ( .A(a1[2]), .ZN(n15) );
  INV_X1 U142 ( .A(n15), .ZN(n16) );
  INV_X1 U143 ( .A(n17), .ZN(n18) );
  INV_X4 U144 ( .A(a2[16]), .ZN(n19) );
  INV_X1 U145 ( .A(n19), .ZN(n20) );
  INV_X2 U146 ( .A(n21), .ZN(n22) );
  INV_X2 U147 ( .A(n23), .ZN(n24) );
  INV_X2 U148 ( .A(n25), .ZN(n26) );
  INV_X2 U149 ( .A(n27), .ZN(n28) );
  INV_X2 U150 ( .A(n29), .ZN(n30) );
  INV_X2 U151 ( .A(n31), .ZN(n32) );
  INV_X2 U152 ( .A(n33), .ZN(n34) );
  INV_X2 U153 ( .A(n35), .ZN(n36) );
  INV_X2 U154 ( .A(n37), .ZN(n38) );
  INV_X2 U155 ( .A(n39), .ZN(n40) );
  INV_X2 U156 ( .A(n41), .ZN(n42) );
  INV_X2 U157 ( .A(n43), .ZN(n44) );
  INV_X2 U158 ( .A(n45), .ZN(n46) );
  INV_X2 U159 ( .A(n47), .ZN(n48) );
  INV_X2 U160 ( .A(n49), .ZN(n50) );
  INV_X2 U161 ( .A(n51), .ZN(n52) );
  INV_X2 U162 ( .A(n53), .ZN(n54) );
  INV_X2 U163 ( .A(n55), .ZN(n56) );
  INV_X2 U164 ( .A(n57), .ZN(n58) );
  INV_X2 U165 ( .A(n59), .ZN(n60) );
  INV_X2 U166 ( .A(n61), .ZN(n62) );
  INV_X2 U167 ( .A(n63), .ZN(n64) );
  INV_X2 U168 ( .A(n65), .ZN(n66) );
  INV_X2 U169 ( .A(n67), .ZN(n68) );
  INV_X2 U170 ( .A(n69), .ZN(n70) );
  INV_X2 U171 ( .A(n71), .ZN(n72) );
  INV_X2 U172 ( .A(n73), .ZN(n74) );
  INV_X2 U173 ( .A(n75), .ZN(n76) );
  INV_X2 U174 ( .A(n77), .ZN(n78) );
  INV_X2 U175 ( .A(n79), .ZN(n80) );
  INV_X2 U176 ( .A(n81), .ZN(n82) );
  INV_X2 U177 ( .A(n83), .ZN(n84) );
  INV_X2 U178 ( .A(n85), .ZN(n86) );
  INV_X2 U179 ( .A(n87), .ZN(n88) );
  INV_X2 U180 ( .A(n89), .ZN(n90) );
  INV_X2 U181 ( .A(n91), .ZN(n92) );
  INV_X2 U182 ( .A(n93), .ZN(n94) );
  INV_X2 U183 ( .A(n95), .ZN(n96) );
  INV_X2 U184 ( .A(n97), .ZN(n98) );
  INV_X2 U185 ( .A(n99), .ZN(n100) );
  INV_X2 U186 ( .A(n101), .ZN(n102) );
  INV_X2 U187 ( .A(n103), .ZN(n104) );
  INV_X2 U188 ( .A(n105), .ZN(n106) );
  INV_X2 U189 ( .A(n107), .ZN(n108) );
  INV_X2 U190 ( .A(n109), .ZN(n110) );
  INV_X2 U191 ( .A(n111), .ZN(n112) );
  INV_X2 U192 ( .A(n113), .ZN(n114) );
  INV_X2 U193 ( .A(n115), .ZN(n116) );
  INV_X2 U194 ( .A(n117), .ZN(n118) );
  INV_X2 U195 ( .A(n119), .ZN(n120) );
  INV_X2 U196 ( .A(n121), .ZN(n122) );
  INV_X2 U197 ( .A(n123), .ZN(n124) );
  INV_X2 U198 ( .A(n125), .ZN(n126) );
  INV_X2 U199 ( .A(n127), .ZN(n128) );
  INV_X2 U200 ( .A(n129), .ZN(n130) );
  INV_X2 U201 ( .A(n131), .ZN(n132) );
  INV_X2 U202 ( .A(n133), .ZN(n134) );
  INV_X2 U203 ( .A(n135), .ZN(n136) );
  INV_X2 U204 ( .A(n137), .ZN(n138) );
  INV_X2 U205 ( .A(n139), .ZN(n140) );
  INV_X2 U206 ( .A(n141), .ZN(n142) );
  INV_X2 U207 ( .A(n143), .ZN(n144) );
  INV_X2 U208 ( .A(n145), .ZN(n146) );
  INV_X2 U209 ( .A(n147), .ZN(n148) );
  INV_X2 U210 ( .A(n149), .ZN(n150) );
  INV_X2 U211 ( .A(n151), .ZN(n152) );
  INV_X2 U212 ( .A(n153), .ZN(n154) );
  INV_X2 U213 ( .A(n155), .ZN(n156) );
  INV_X2 U214 ( .A(n157), .ZN(n158) );
  INV_X2 U215 ( .A(n159), .ZN(n160) );
  INV_X2 U216 ( .A(n161), .ZN(n162) );
  INV_X2 U217 ( .A(n163), .ZN(n164) );
  INV_X2 U218 ( .A(n165), .ZN(n166) );
  INV_X2 U219 ( .A(n167), .ZN(n168) );
  INV_X2 U220 ( .A(n169), .ZN(n170) );
  INV_X2 U221 ( .A(n171), .ZN(n172) );
  INV_X2 U222 ( .A(n173), .ZN(n174) );
  INV_X2 U223 ( .A(n175), .ZN(n176) );
  INV_X2 U224 ( .A(n177), .ZN(n178) );
  INV_X2 U225 ( .A(n179), .ZN(n180) );
  INV_X2 U226 ( .A(n181), .ZN(n182) );
  INV_X2 U227 ( .A(n183), .ZN(n184) );
  INV_X2 U228 ( .A(n185), .ZN(n186) );
  INV_X2 U229 ( .A(n187), .ZN(n188) );
  INV_X2 U230 ( .A(n189), .ZN(n190) );
  INV_X2 U231 ( .A(n191), .ZN(n192) );
  INV_X2 U232 ( .A(n193), .ZN(n194) );
  INV_X2 U233 ( .A(n195), .ZN(n196) );
  INV_X2 U234 ( .A(n197), .ZN(n198) );
  INV_X2 U235 ( .A(n199), .ZN(n200) );
  INV_X2 U236 ( .A(n201), .ZN(n202) );
  INV_X2 U237 ( .A(n203), .ZN(n204) );
  INV_X2 U238 ( .A(n205), .ZN(n206) );
  INV_X2 U239 ( .A(n207), .ZN(n208) );
  INV_X2 U240 ( .A(n209), .ZN(n210) );
  INV_X2 U241 ( .A(n211), .ZN(n212) );
  INV_X2 U242 ( .A(n213), .ZN(n214) );
  INV_X2 U243 ( .A(n215), .ZN(n216) );
  INV_X2 U244 ( .A(n217), .ZN(n218) );
  INV_X2 U245 ( .A(n219), .ZN(n220) );
  INV_X2 U246 ( .A(n221), .ZN(n222) );
  INV_X2 U247 ( .A(n223), .ZN(n224) );
  INV_X2 U248 ( .A(n225), .ZN(n226) );
  INV_X2 U249 ( .A(n227), .ZN(n228) );
  INV_X2 U250 ( .A(n229), .ZN(n230) );
  INV_X2 U251 ( .A(n231), .ZN(n232) );
  INV_X2 U252 ( .A(n233), .ZN(n234) );
  INV_X2 U253 ( .A(n235), .ZN(n236) );
  INV_X2 U254 ( .A(n237), .ZN(n238) );
  INV_X2 U255 ( .A(n239), .ZN(n240) );
  INV_X2 U256 ( .A(n241), .ZN(n242) );
  INV_X2 U257 ( .A(n243), .ZN(n244) );
  INV_X2 U258 ( .A(n245), .ZN(n246) );
  INV_X2 U259 ( .A(n247), .ZN(n248) );
  INV_X2 U260 ( .A(n249), .ZN(n250) );
  INV_X2 U261 ( .A(n251), .ZN(n252) );
  INV_X2 U262 ( .A(n253), .ZN(n254) );
  INV_X2 U263 ( .A(n255), .ZN(n256) );
  INV_X2 U264 ( .A(n257), .ZN(n258) );
  INV_X2 U265 ( .A(n259), .ZN(n260) );
  INV_X2 U266 ( .A(n261), .ZN(n262) );
  INV_X2 U267 ( .A(n263), .ZN(n264) );
  INV_X2 U268 ( .A(n265), .ZN(n266) );
  INV_X2 U269 ( .A(n267), .ZN(n268) );
endmodule

