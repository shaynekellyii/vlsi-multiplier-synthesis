
module mul32_3_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n262, n265, n268, n271, n274, n277, n280, n283, n286, n289, n291,
         n293, n295, n297, n299, n307, n313, n315, n317, n319, n321, n323,
         n325, n327, n329, n331, n333, n336, n339, n342, n345, n348, n351,
         n354, n357, n360, n363, n366, n368, n370, n372, n374, n376, n378,
         n380, n382, n384, n386, n388, n390, n393, n397, n400, n403, n406,
         n409, n412, n415, n418, n421, n424, n427, n430, n433, n436, n439,
         n442, n445, n448, n451, n454, n457, n460, n463, n466, n469, n472,
         n475, n478, n481, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n552, n553, n554, n555, n556, n557, n558,
         n560, n561, n562, n563, n564, n565, n566, n568, n569, n570, n571,
         n572, n573, n574, n576, n577, n578, n579, n580, n581, n582, n584,
         n585, n586, n587, n588, n589, n590, n592, n593, n594, n595, n596,
         n597, n598, n600, n601, n602, n603, n604, n605, n606, n608, n609,
         n610, n611, n612, n613, n614, n616, n617, n618, n619, n620, n621,
         n622, n624, n625, n626, n627, n628, n629, n630, n632, n633, n634,
         n635, n636, n637, n638, n640, n641, n642, n643, n644, n645, n646,
         n648, n649, n650, n651, n652, n653, n654, n656, n657, n658, n659,
         n660, n661, n662, n664, n665, n666, n667, n668, n669, n670, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1376, n1377, n1379, n1380,
         n1382, n1383, n1385, n1386, n1388, n1389, n1391, n1392, n1394, n1395,
         n1397, n1398, n1400, n1401, n1403, n1404, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1518, n1519, n1520, n1521, n1522, n1523, n1526,
         n1527, n1528, n1529, n1530, n1531, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1564,
         n1565, n1568, n1569, n1570, n1571, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1584, n1585, n1586, n1587, n1588, n1589, n1592,
         n1593, n1594, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1620, n1621, n1622, n1623, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1635, n1636, n1637, n1638, n1639,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237;
  assign n262 = a[2];
  assign n265 = a[5];
  assign n268 = a[8];
  assign n271 = a[11];
  assign n274 = a[14];
  assign n277 = a[17];
  assign n280 = a[20];
  assign n283 = a[23];
  assign n286 = a[26];
  assign n289 = a[29];
  assign n390 = b[0];
  assign n393 = b[1];
  assign n397 = b[2];
  assign n400 = b[3];
  assign n403 = b[4];
  assign n406 = b[5];
  assign n409 = b[6];
  assign n412 = b[7];
  assign n415 = b[8];
  assign n418 = b[9];
  assign n421 = b[10];
  assign n424 = b[11];
  assign n427 = b[12];
  assign n430 = b[13];
  assign n433 = b[14];
  assign n436 = b[15];
  assign n439 = b[16];
  assign n442 = b[17];
  assign n445 = b[18];
  assign n448 = b[19];
  assign n451 = b[20];
  assign n454 = b[21];
  assign n457 = b[22];
  assign n460 = b[23];
  assign n463 = b[24];
  assign n466 = b[25];
  assign n469 = b[26];
  assign n472 = b[27];
  assign n475 = b[28];
  assign n478 = b[29];
  assign n481 = b[30];
  assign n484 = b[31];

  XOR2_X2 U304 ( .A(n717), .B(n716), .Z(n485) );
  FA_X1 U305 ( .A(n719), .B(n718), .CI(n520), .CO(n519), .S(product[62]) );
  FA_X1 U306 ( .A(n720), .B(n721), .CI(n521), .CO(n520), .S(product[61]) );
  FA_X1 U307 ( .A(n725), .B(n722), .CI(n522), .CO(n521), .S(product[60]) );
  FA_X1 U308 ( .A(n726), .B(n728), .CI(n523), .CO(n522), .S(product[59]) );
  FA_X1 U313 ( .A(n743), .B(n739), .CI(n526), .CO(n525), .S(product[56]) );
  FA_X1 U314 ( .A(n744), .B(n749), .CI(n527), .CO(n526), .S(product[55]) );
  FA_X1 U315 ( .A(n750), .B(n757), .CI(n528), .CO(n527), .S(product[54]) );
  FA_X1 U316 ( .A(n758), .B(n764), .CI(n529), .CO(n528), .S(product[53]) );
  FA_X1 U319 ( .A(n783), .B(n791), .CI(n532), .CO(n531), .S(product[50]) );
  FA_X1 U320 ( .A(n792), .B(n801), .CI(n533), .CO(n532), .S(product[49]) );
  FA_X1 U323 ( .A(n825), .B(n836), .CI(n536), .CO(n535), .S(product[46]) );
  FA_X1 U324 ( .A(n837), .B(n850), .CI(n537), .CO(n536), .S(product[45]) );
  FA_X1 U325 ( .A(n851), .B(n863), .CI(n538), .CO(n537), .S(product[44]) );
  FA_X1 U326 ( .A(n864), .B(n877), .CI(n539), .CO(n538), .S(product[43]) );
  FA_X1 U327 ( .A(n878), .B(n893), .CI(n540), .CO(n539), .S(product[42]) );
  FA_X1 U328 ( .A(n894), .B(n909), .CI(n541), .CO(n540), .S(product[41]) );
  FA_X1 U333 ( .A(n979), .B(n996), .CI(n546), .CO(n545), .S(product[36]) );
  FA_X1 U334 ( .A(n997), .B(n1014), .CI(n547), .CO(n546), .S(product[35]) );
  NAND2_X4 U337 ( .A1(n683), .A2(n549), .ZN(n486) );
  NOR2_X4 U339 ( .A1(n1015), .A2(n1032), .ZN(n548) );
  NAND2_X4 U340 ( .A1(n1015), .A2(n1032), .ZN(n549) );
  NAND2_X4 U345 ( .A1(n684), .A2(n554), .ZN(n487) );
  NOR2_X4 U347 ( .A1(n1033), .A2(n1050), .ZN(n553) );
  NAND2_X4 U348 ( .A1(n1033), .A2(n1050), .ZN(n554) );
  NAND2_X4 U351 ( .A1(n685), .A2(n557), .ZN(n488) );
  NOR2_X4 U353 ( .A1(n1051), .A2(n1068), .ZN(n556) );
  NAND2_X4 U354 ( .A1(n1051), .A2(n1068), .ZN(n557) );
  AOI21_X4 U356 ( .B1(n563), .B2(n686), .A(n560), .ZN(n558) );
  NAND2_X4 U359 ( .A1(n686), .A2(n562), .ZN(n489) );
  NOR2_X4 U361 ( .A1(n1069), .A2(n1086), .ZN(n561) );
  NAND2_X4 U362 ( .A1(n1069), .A2(n1086), .ZN(n562) );
  NAND2_X4 U365 ( .A1(n687), .A2(n565), .ZN(n490) );
  NOR2_X4 U367 ( .A1(n1087), .A2(n1104), .ZN(n564) );
  NAND2_X4 U368 ( .A1(n1087), .A2(n1104), .ZN(n565) );
  NAND2_X4 U373 ( .A1(n688), .A2(n570), .ZN(n491) );
  NOR2_X4 U375 ( .A1(n1105), .A2(n1122), .ZN(n569) );
  NAND2_X4 U376 ( .A1(n1105), .A2(n1122), .ZN(n570) );
  NAND2_X4 U379 ( .A1(n689), .A2(n573), .ZN(n492) );
  NOR2_X4 U381 ( .A1(n1123), .A2(n1140), .ZN(n572) );
  NAND2_X4 U382 ( .A1(n1123), .A2(n1140), .ZN(n573) );
  NAND2_X4 U387 ( .A1(n690), .A2(n578), .ZN(n493) );
  NOR2_X4 U389 ( .A1(n1141), .A2(n1158), .ZN(n577) );
  NAND2_X4 U390 ( .A1(n1141), .A2(n1158), .ZN(n578) );
  NAND2_X4 U393 ( .A1(n691), .A2(n581), .ZN(n494) );
  NOR2_X4 U395 ( .A1(n1159), .A2(n1174), .ZN(n580) );
  NAND2_X4 U396 ( .A1(n1159), .A2(n1174), .ZN(n581) );
  AOI21_X4 U398 ( .B1(n587), .B2(n692), .A(n584), .ZN(n582) );
  NAND2_X4 U401 ( .A1(n692), .A2(n586), .ZN(n495) );
  NOR2_X4 U403 ( .A1(n1175), .A2(n1190), .ZN(n585) );
  NAND2_X4 U404 ( .A1(n1175), .A2(n1190), .ZN(n586) );
  NAND2_X4 U407 ( .A1(n693), .A2(n589), .ZN(n496) );
  NOR2_X4 U409 ( .A1(n1191), .A2(n1206), .ZN(n588) );
  NAND2_X4 U412 ( .A1(n1191), .A2(n1206), .ZN(n589) );
  NAND2_X4 U417 ( .A1(n694), .A2(n594), .ZN(n497) );
  NOR2_X4 U419 ( .A1(n1207), .A2(n1220), .ZN(n593) );
  NAND2_X4 U420 ( .A1(n1207), .A2(n1220), .ZN(n594) );
  NAND2_X4 U423 ( .A1(n695), .A2(n597), .ZN(n498) );
  NOR2_X4 U425 ( .A1(n1221), .A2(n1234), .ZN(n596) );
  NAND2_X4 U426 ( .A1(n1221), .A2(n1234), .ZN(n597) );
  NAND2_X4 U431 ( .A1(n696), .A2(n602), .ZN(n499) );
  NOR2_X4 U433 ( .A1(n1235), .A2(n1248), .ZN(n601) );
  NAND2_X4 U434 ( .A1(n1235), .A2(n1248), .ZN(n602) );
  XOR2_X2 U435 ( .A(n606), .B(n500), .Z(product[20]) );
  NAND2_X4 U437 ( .A1(n697), .A2(n605), .ZN(n500) );
  NOR2_X4 U439 ( .A1(n1249), .A2(n1260), .ZN(n604) );
  NAND2_X4 U440 ( .A1(n1249), .A2(n1260), .ZN(n605) );
  AOI21_X4 U442 ( .B1(n611), .B2(n698), .A(n608), .ZN(n606) );
  NAND2_X4 U445 ( .A1(n698), .A2(n610), .ZN(n501) );
  NOR2_X4 U447 ( .A1(n1261), .A2(n1272), .ZN(n609) );
  NAND2_X4 U448 ( .A1(n1261), .A2(n1272), .ZN(n610) );
  NAND2_X4 U451 ( .A1(n699), .A2(n613), .ZN(n502) );
  NOR2_X4 U453 ( .A1(n1273), .A2(n1284), .ZN(n612) );
  NAND2_X4 U454 ( .A1(n1273), .A2(n1284), .ZN(n613) );
  AOI21_X4 U456 ( .B1(n619), .B2(n700), .A(n616), .ZN(n614) );
  NAND2_X4 U459 ( .A1(n700), .A2(n618), .ZN(n503) );
  NOR2_X4 U461 ( .A1(n1285), .A2(n1294), .ZN(n617) );
  NAND2_X4 U462 ( .A1(n1285), .A2(n1294), .ZN(n618) );
  NAND2_X4 U465 ( .A1(n701), .A2(n621), .ZN(n504) );
  NOR2_X4 U467 ( .A1(n1295), .A2(n1304), .ZN(n620) );
  NAND2_X4 U468 ( .A1(n1295), .A2(n1304), .ZN(n621) );
  AOI21_X4 U470 ( .B1(n627), .B2(n702), .A(n624), .ZN(n622) );
  NAND2_X4 U473 ( .A1(n702), .A2(n626), .ZN(n505) );
  NOR2_X4 U475 ( .A1(n1305), .A2(n1314), .ZN(n625) );
  NAND2_X4 U476 ( .A1(n1305), .A2(n1314), .ZN(n626) );
  NAND2_X4 U479 ( .A1(n703), .A2(n629), .ZN(n506) );
  NOR2_X4 U481 ( .A1(n1315), .A2(n1322), .ZN(n628) );
  NAND2_X4 U482 ( .A1(n1315), .A2(n1322), .ZN(n629) );
  AOI21_X4 U484 ( .B1(n635), .B2(n704), .A(n632), .ZN(n630) );
  NAND2_X4 U487 ( .A1(n704), .A2(n634), .ZN(n507) );
  XOR2_X2 U491 ( .A(n638), .B(n508), .Z(product[12]) );
  NAND2_X4 U493 ( .A1(n705), .A2(n637), .ZN(n508) );
  NOR2_X4 U495 ( .A1(n1331), .A2(n1338), .ZN(n636) );
  NAND2_X4 U496 ( .A1(n1331), .A2(n1338), .ZN(n637) );
  AOI21_X4 U498 ( .B1(n643), .B2(n706), .A(n640), .ZN(n638) );
  NAND2_X4 U501 ( .A1(n706), .A2(n642), .ZN(n509) );
  NOR2_X4 U503 ( .A1(n1339), .A2(n1344), .ZN(n641) );
  NAND2_X4 U504 ( .A1(n1339), .A2(n1344), .ZN(n642) );
  NAND2_X4 U507 ( .A1(n707), .A2(n645), .ZN(n510) );
  NOR2_X4 U509 ( .A1(n1345), .A2(n1350), .ZN(n644) );
  NAND2_X4 U510 ( .A1(n1345), .A2(n1350), .ZN(n645) );
  NAND2_X4 U515 ( .A1(n708), .A2(n650), .ZN(n511) );
  NAND2_X4 U518 ( .A1(n1351), .A2(n1356), .ZN(n650) );
  XOR2_X2 U519 ( .A(n654), .B(n512), .Z(product[8]) );
  NAND2_X4 U521 ( .A1(n709), .A2(n653), .ZN(n512) );
  NOR2_X4 U523 ( .A1(n1357), .A2(n1360), .ZN(n652) );
  NAND2_X4 U524 ( .A1(n1357), .A2(n1360), .ZN(n653) );
  XNOR2_X2 U525 ( .A(n513), .B(n659), .ZN(product[7]) );
  AOI21_X4 U526 ( .B1(n710), .B2(n659), .A(n656), .ZN(n654) );
  NAND2_X4 U529 ( .A1(n710), .A2(n658), .ZN(n513) );
  NOR2_X4 U531 ( .A1(n1361), .A2(n1364), .ZN(n657) );
  NAND2_X4 U532 ( .A1(n1361), .A2(n1364), .ZN(n658) );
  XOR2_X2 U533 ( .A(n514), .B(n662), .Z(product[6]) );
  NAND2_X4 U535 ( .A1(n711), .A2(n661), .ZN(n514) );
  NOR2_X4 U537 ( .A1(n1365), .A2(n2087), .ZN(n660) );
  NAND2_X4 U538 ( .A1(n1365), .A2(n2087), .ZN(n661) );
  XNOR2_X2 U539 ( .A(n515), .B(n667), .ZN(product[5]) );
  AOI21_X4 U540 ( .B1(n712), .B2(n667), .A(n664), .ZN(n662) );
  NAND2_X4 U543 ( .A1(n712), .A2(n666), .ZN(n515) );
  NOR2_X4 U545 ( .A1(n2088), .A2(n1369), .ZN(n665) );
  NAND2_X4 U546 ( .A1(n2088), .A2(n1369), .ZN(n666) );
  XOR2_X2 U547 ( .A(n516), .B(n670), .Z(product[4]) );
  OAI21_X4 U548 ( .B1(n670), .B2(n668), .A(n669), .ZN(n667) );
  NAND2_X4 U549 ( .A1(n713), .A2(n669), .ZN(n516) );
  NOR2_X4 U551 ( .A1(n1371), .A2(n2089), .ZN(n668) );
  NAND2_X4 U552 ( .A1(n1371), .A2(n2089), .ZN(n669) );
  XNOR2_X2 U553 ( .A(n517), .B(n675), .ZN(product[3]) );
  AOI21_X4 U554 ( .B1(n675), .B2(n714), .A(n672), .ZN(n670) );
  NAND2_X4 U557 ( .A1(n714), .A2(n674), .ZN(n517) );
  NOR2_X4 U559 ( .A1(n2090), .A2(n1373), .ZN(n673) );
  NAND2_X4 U560 ( .A1(n2090), .A2(n1373), .ZN(n674) );
  XOR2_X2 U561 ( .A(n676), .B(n677), .Z(product[2]) );
  NOR2_X4 U562 ( .A1(n676), .A2(n677), .ZN(n675) );
  XNOR2_X2 U564 ( .A(n679), .B(n680), .ZN(product[1]) );
  NAND2_X4 U565 ( .A1(n678), .A2(n680), .ZN(n677) );
  NAND2_X4 U570 ( .A1(n715), .A2(n682), .ZN(n518) );
  NOR2_X4 U572 ( .A1(n2093), .A2(n262), .ZN(n681) );
  FA_X1 U576 ( .A(n1721), .B(n1745), .CI(n723), .CO(n719), .S(n720) );
  FA_X1 U577 ( .A(n727), .B(n1722), .CI(n1746), .CO(n721), .S(n722) );
  FA_X1 U579 ( .A(n1747), .B(n727), .CI(n730), .CO(n725), .S(n726) );
  FA_X1 U581 ( .A(n734), .B(n1748), .CI(n731), .CO(n728), .S(n729) );
  FA_X1 U582 ( .A(n736), .B(n1779), .CI(n1723), .CO(n730), .S(n731) );
  FA_X1 U583 ( .A(n740), .B(n1749), .CI(n735), .CO(n732), .S(n733) );
  FA_X1 U584 ( .A(n742), .B(n1724), .CI(n1780), .CO(n734), .S(n735) );
  FA_X1 U586 ( .A(n741), .B(n747), .CI(n745), .CO(n738), .S(n739) );
  FA_X1 U587 ( .A(n1781), .B(n742), .CI(n1750), .CO(n740), .S(n741) );
  FA_X1 U589 ( .A(n751), .B(n748), .CI(n746), .CO(n743), .S(n744) );
  FA_X1 U590 ( .A(n1751), .B(n1782), .CI(n753), .CO(n745), .S(n746) );
  FA_X1 U591 ( .A(n755), .B(n1814), .CI(n1725), .CO(n747), .S(n748) );
  FA_X1 U592 ( .A(n759), .B(n754), .CI(n752), .CO(n749), .S(n750) );
  FA_X1 U593 ( .A(n1752), .B(n1783), .CI(n761), .CO(n751), .S(n752) );
  FA_X1 U594 ( .A(n763), .B(n1726), .CI(n1815), .CO(n753), .S(n754) );
  FA_X1 U596 ( .A(n766), .B(n762), .CI(n760), .CO(n757), .S(n758) );
  FA_X1 U597 ( .A(n770), .B(n1753), .CI(n768), .CO(n759), .S(n760) );
  FA_X1 U598 ( .A(n1816), .B(n763), .CI(n1784), .CO(n761), .S(n762) );
  FA_X1 U600 ( .A(n774), .B(n769), .CI(n767), .CO(n764), .S(n765) );
  FA_X1 U601 ( .A(n771), .B(n778), .CI(n776), .CO(n766), .S(n767) );
  FA_X1 U602 ( .A(n1785), .B(n1754), .CI(n1817), .CO(n768), .S(n769) );
  FA_X1 U603 ( .A(n780), .B(n1849), .CI(n1727), .CO(n770), .S(n771) );
  FA_X1 U604 ( .A(n784), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U605 ( .A(n779), .B(n788), .CI(n786), .CO(n774), .S(n775) );
  FA_X1 U606 ( .A(n1786), .B(n1755), .CI(n1818), .CO(n776), .S(n777) );
  FA_X1 U607 ( .A(n790), .B(n1728), .CI(n1850), .CO(n778), .S(n779) );
  FA_X1 U609 ( .A(n793), .B(n787), .CI(n785), .CO(n782), .S(n783) );
  FA_X1 U610 ( .A(n789), .B(n797), .CI(n795), .CO(n784), .S(n785) );
  FA_X1 U611 ( .A(n1787), .B(n1819), .CI(n799), .CO(n786), .S(n787) );
  FA_X1 U612 ( .A(n1851), .B(n790), .CI(n1756), .CO(n788), .S(n789) );
  FA_X1 U614 ( .A(n803), .B(n796), .CI(n794), .CO(n791), .S(n792) );
  FA_X1 U615 ( .A(n798), .B(n807), .CI(n805), .CO(n793), .S(n794) );
  FA_X1 U616 ( .A(n809), .B(n1820), .CI(n800), .CO(n795), .S(n796) );
  FA_X1 U617 ( .A(n1852), .B(n1757), .CI(n1788), .CO(n797), .S(n798) );
  FA_X1 U618 ( .A(n811), .B(n1884), .CI(n1729), .CO(n799), .S(n800) );
  FA_X1 U619 ( .A(n815), .B(n806), .CI(n804), .CO(n801), .S(n802) );
  FA_X1 U620 ( .A(n808), .B(n819), .CI(n817), .CO(n803), .S(n804) );
  FA_X1 U621 ( .A(n821), .B(n1758), .CI(n810), .CO(n805), .S(n806) );
  FA_X1 U622 ( .A(n1853), .B(n1789), .CI(n1821), .CO(n807), .S(n808) );
  FA_X1 U623 ( .A(n823), .B(n1730), .CI(n1885), .CO(n809), .S(n810) );
  FA_X1 U625 ( .A(n826), .B(n818), .CI(n816), .CO(n813), .S(n814) );
  FA_X1 U626 ( .A(n820), .B(n822), .CI(n828), .CO(n815), .S(n816) );
  FA_X1 U627 ( .A(n832), .B(n1759), .CI(n830), .CO(n817), .S(n818) );
  FA_X1 U628 ( .A(n1822), .B(n1790), .CI(n1854), .CO(n819), .S(n820) );
  FA_X1 U629 ( .A(n834), .B(n823), .CI(n1886), .CO(n821), .S(n822) );
  FA_X1 U631 ( .A(n838), .B(n829), .CI(n827), .CO(n824), .S(n825) );
  FA_X1 U632 ( .A(n842), .B(n833), .CI(n840), .CO(n826), .S(n827) );
  FA_X1 U633 ( .A(n844), .B(n846), .CI(n831), .CO(n828), .S(n829) );
  FA_X1 U634 ( .A(n1823), .B(n1760), .CI(n1887), .CO(n830), .S(n831) );
  FA_X1 U635 ( .A(n1855), .B(n1791), .CI(n835), .CO(n832), .S(n833) );
  FA_X1 U636 ( .A(n848), .B(n1919), .CI(n1731), .CO(n834), .S(n835) );
  FA_X1 U637 ( .A(n852), .B(n841), .CI(n839), .CO(n836), .S(n837) );
  FA_X1 U638 ( .A(n843), .B(n856), .CI(n854), .CO(n838), .S(n839) );
  FA_X1 U639 ( .A(n858), .B(n847), .CI(n845), .CO(n840), .S(n841) );
  FA_X1 U640 ( .A(n1761), .B(n1824), .CI(n860), .CO(n842), .S(n843) );
  FA_X1 U641 ( .A(n1888), .B(n1792), .CI(n1856), .CO(n844), .S(n845) );
  FA_X1 U642 ( .A(n1732), .B(n862), .CI(n1920), .CO(n846), .S(n847) );
  FA_X1 U644 ( .A(n865), .B(n855), .CI(n853), .CO(n850), .S(n851) );
  FA_X1 U645 ( .A(n857), .B(n869), .CI(n867), .CO(n852), .S(n853) );
  FA_X1 U646 ( .A(n861), .B(n871), .CI(n859), .CO(n854), .S(n855) );
  FA_X1 U647 ( .A(n1857), .B(n1762), .CI(n873), .CO(n856), .S(n857) );
  FA_X1 U648 ( .A(n1889), .B(n1793), .CI(n875), .CO(n858), .S(n859) );
  FA_X1 U649 ( .A(n1921), .B(n862), .CI(n1825), .CO(n860), .S(n861) );
  FA_X1 U651 ( .A(n879), .B(n868), .CI(n866), .CO(n863), .S(n864) );
  FA_X1 U652 ( .A(n870), .B(n883), .CI(n881), .CO(n865), .S(n866) );
  FA_X1 U653 ( .A(n874), .B(n885), .CI(n872), .CO(n867), .S(n868) );
  FA_X1 U654 ( .A(n889), .B(n876), .CI(n887), .CO(n869), .S(n870) );
  FA_X1 U655 ( .A(n1858), .B(n1922), .CI(n1890), .CO(n871), .S(n872) );
  FA_X1 U656 ( .A(n1826), .B(n1763), .CI(n1794), .CO(n873), .S(n874) );
  FA_X1 U657 ( .A(n891), .B(n3208), .CI(n1733), .CO(n875), .S(n876) );
  FA_X1 U658 ( .A(n895), .B(n882), .CI(n880), .CO(n877), .S(n878) );
  FA_X1 U659 ( .A(n884), .B(n899), .CI(n897), .CO(n879), .S(n880) );
  FA_X1 U660 ( .A(n888), .B(n901), .CI(n886), .CO(n881), .S(n882) );
  FA_X1 U661 ( .A(n890), .B(n905), .CI(n903), .CO(n883), .S(n884) );
  FA_X1 U662 ( .A(n1891), .B(n1859), .CI(n1923), .CO(n885), .S(n886) );
  FA_X1 U663 ( .A(n1827), .B(n1764), .CI(n1795), .CO(n887), .S(n888) );
  FA_X1 U664 ( .A(n907), .B(n892), .CI(n1955), .CO(n889), .S(n890) );
  FA_X1 U666 ( .A(n911), .B(n898), .CI(n896), .CO(n893), .S(n894) );
  FA_X1 U667 ( .A(n900), .B(n915), .CI(n913), .CO(n895), .S(n896) );
  FA_X1 U668 ( .A(n904), .B(n917), .CI(n902), .CO(n897), .S(n898) );
  FA_X1 U669 ( .A(n921), .B(n906), .CI(n919), .CO(n899), .S(n900) );
  FA_X1 U670 ( .A(n1892), .B(n1796), .CI(n1924), .CO(n901), .S(n902) );
  FA_X1 U671 ( .A(n1828), .B(n1956), .CI(n1860), .CO(n903), .S(n904) );
  FA_X1 U672 ( .A(n908), .B(n1734), .CI(n923), .CO(n905), .S(n906) );
  FA_X1 U674 ( .A(n927), .B(n914), .CI(n912), .CO(n909), .S(n910) );
  FA_X1 U675 ( .A(n916), .B(n931), .CI(n929), .CO(n911), .S(n912) );
  FA_X1 U676 ( .A(n920), .B(n933), .CI(n918), .CO(n913), .S(n914) );
  FA_X1 U677 ( .A(n935), .B(n937), .CI(n922), .CO(n915), .S(n916) );
  FA_X1 U678 ( .A(n1893), .B(n1829), .CI(n1957), .CO(n917), .S(n918) );
  FA_X1 U679 ( .A(n1925), .B(n1861), .CI(n939), .CO(n919), .S(n920) );
  FA_X1 U680 ( .A(n1765), .B(n1797), .CI(n924), .CO(n921), .S(n922) );
  FA_X1 U681 ( .A(n941), .B(n3216), .CI(n1735), .CO(n923), .S(n924) );
  FA_X1 U682 ( .A(n945), .B(n930), .CI(n928), .CO(n925), .S(n926) );
  FA_X1 U683 ( .A(n932), .B(n949), .CI(n947), .CO(n927), .S(n928) );
  FA_X1 U684 ( .A(n951), .B(n936), .CI(n934), .CO(n929), .S(n930) );
  FA_X1 U685 ( .A(n953), .B(n955), .CI(n938), .CO(n931), .S(n932) );
  FA_X1 U686 ( .A(n957), .B(n1894), .CI(n940), .CO(n933), .S(n934) );
  FA_X1 U687 ( .A(n1926), .B(n1830), .CI(n1958), .CO(n935), .S(n936) );
  FA_X1 U688 ( .A(n1798), .B(n1990), .CI(n1862), .CO(n937), .S(n938) );
  FA_X1 U689 ( .A(n1736), .B(n959), .CI(n1766), .CO(n939), .S(n940) );
  FA_X1 U691 ( .A(n962), .B(n948), .CI(n946), .CO(n943), .S(n944) );
  FA_X1 U692 ( .A(n950), .B(n966), .CI(n964), .CO(n945), .S(n946) );
  FA_X1 U693 ( .A(n968), .B(n954), .CI(n952), .CO(n947), .S(n948) );
  FA_X1 U694 ( .A(n970), .B(n972), .CI(n956), .CO(n949), .S(n950) );
  FA_X1 U695 ( .A(n974), .B(n1895), .CI(n958), .CO(n951), .S(n952) );
  FA_X1 U696 ( .A(n1927), .B(n1831), .CI(n1959), .CO(n953), .S(n954) );
  FA_X1 U697 ( .A(n1767), .B(n1991), .CI(n1863), .CO(n955), .S(n956) );
  FA_X1 U698 ( .A(n1799), .B(n959), .CI(n976), .CO(n957), .S(n958) );
  FA_X1 U700 ( .A(n980), .B(n965), .CI(n963), .CO(n960), .S(n961) );
  FA_X1 U701 ( .A(n967), .B(n969), .CI(n982), .CO(n962), .S(n963) );
  FA_X1 U702 ( .A(n986), .B(n971), .CI(n984), .CO(n964), .S(n965) );
  FA_X1 U703 ( .A(n975), .B(n988), .CI(n973), .CO(n966), .S(n967) );
  FA_X1 U704 ( .A(n992), .B(n1960), .CI(n990), .CO(n968), .S(n969) );
  FA_X1 U705 ( .A(n1928), .B(n1992), .CI(n994), .CO(n970), .S(n971) );
  FA_X1 U706 ( .A(n1896), .B(n977), .CI(n1864), .CO(n972), .S(n973) );
  FA_X1 U707 ( .A(n1832), .B(n1768), .CI(n1800), .CO(n974), .S(n975) );
  FA_X1 U708 ( .A(n2024), .B(n3209), .CI(n1737), .CO(n976), .S(n977) );
  FA_X1 U709 ( .A(n998), .B(n983), .CI(n981), .CO(n978), .S(n979) );
  FA_X1 U710 ( .A(n985), .B(n987), .CI(n1000), .CO(n980), .S(n981) );
  FA_X1 U711 ( .A(n1004), .B(n989), .CI(n1002), .CO(n982), .S(n983) );
  FA_X1 U712 ( .A(n993), .B(n1006), .CI(n991), .CO(n984), .S(n985) );
  FA_X1 U713 ( .A(n1010), .B(n995), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U714 ( .A(n1865), .B(n1929), .CI(n1961), .CO(n988), .S(n989) );
  FA_X1 U715 ( .A(n1897), .B(n1012), .CI(n1993), .CO(n990), .S(n991) );
  FA_X1 U716 ( .A(n2025), .B(n1769), .CI(n1833), .CO(n992), .S(n993) );
  FA_X1 U717 ( .A(n1738), .B(n262), .CI(n1801), .CO(n994), .S(n995) );
  FA_X1 U718 ( .A(n1016), .B(n1001), .CI(n999), .CO(n996), .S(n997) );
  FA_X1 U719 ( .A(n1003), .B(n1005), .CI(n1018), .CO(n998), .S(n999) );
  FA_X1 U720 ( .A(n1022), .B(n1009), .CI(n1020), .CO(n1000), .S(n1001) );
  FA_X1 U721 ( .A(n1011), .B(n1024), .CI(n1007), .CO(n1002), .S(n1003) );
  FA_X1 U722 ( .A(n1028), .B(n1013), .CI(n1026), .CO(n1004), .S(n1005) );
  FA_X1 U723 ( .A(n1866), .B(n1930), .CI(n1962), .CO(n1006), .S(n1007) );
  FA_X1 U724 ( .A(n1994), .B(n1898), .CI(n1030), .CO(n1008), .S(n1009) );
  FA_X1 U725 ( .A(n2026), .B(n1834), .CI(n1802), .CO(n1010), .S(n1011) );
  FA_X1 U726 ( .A(n1739), .B(n262), .CI(n1770), .CO(n1012), .S(n1013) );
  FA_X1 U727 ( .A(n1034), .B(n1019), .CI(n1017), .CO(n1014), .S(n1015) );
  FA_X1 U728 ( .A(n1021), .B(n1023), .CI(n1036), .CO(n1016), .S(n1017) );
  FA_X1 U729 ( .A(n1040), .B(n1027), .CI(n1038), .CO(n1018), .S(n1019) );
  FA_X1 U730 ( .A(n1029), .B(n1042), .CI(n1025), .CO(n1020), .S(n1021) );
  FA_X1 U731 ( .A(n1046), .B(n1031), .CI(n1044), .CO(n1022), .S(n1023) );
  FA_X1 U732 ( .A(n1963), .B(n1899), .CI(n1995), .CO(n1024), .S(n1025) );
  FA_X1 U733 ( .A(n2027), .B(n1931), .CI(n1048), .CO(n1026), .S(n1027) );
  FA_X1 U734 ( .A(n1867), .B(n1803), .CI(n1835), .CO(n1028), .S(n1029) );
  FA_X1 U735 ( .A(n1740), .B(n262), .CI(n1771), .CO(n1030), .S(n1031) );
  FA_X1 U736 ( .A(n1052), .B(n1037), .CI(n1035), .CO(n1032), .S(n1033) );
  FA_X1 U737 ( .A(n1039), .B(n1041), .CI(n1054), .CO(n1034), .S(n1035) );
  FA_X1 U738 ( .A(n1058), .B(n1045), .CI(n1056), .CO(n1036), .S(n1037) );
  FA_X1 U739 ( .A(n1047), .B(n1060), .CI(n1043), .CO(n1038), .S(n1039) );
  FA_X1 U740 ( .A(n1064), .B(n1049), .CI(n1062), .CO(n1040), .S(n1041) );
  FA_X1 U741 ( .A(n1900), .B(n1964), .CI(n1066), .CO(n1042), .S(n1043) );
  FA_X1 U742 ( .A(n2028), .B(n1932), .CI(n1996), .CO(n1044), .S(n1045) );
  FA_X1 U743 ( .A(n2060), .B(n1836), .CI(n1868), .CO(n1046), .S(n1047) );
  FA_X1 U744 ( .A(n1772), .B(n1741), .CI(n1804), .CO(n1048), .S(n1049) );
  FA_X1 U745 ( .A(n1070), .B(n1055), .CI(n1053), .CO(n1050), .S(n1051) );
  FA_X1 U746 ( .A(n1057), .B(n1059), .CI(n1072), .CO(n1052), .S(n1053) );
  FA_X1 U747 ( .A(n1076), .B(n1063), .CI(n1074), .CO(n1054), .S(n1055) );
  FA_X1 U748 ( .A(n1065), .B(n1078), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U749 ( .A(n1067), .B(n1082), .CI(n1080), .CO(n1058), .S(n1059) );
  FA_X1 U750 ( .A(n1933), .B(n1965), .CI(n1997), .CO(n1060), .S(n1061) );
  FA_X1 U751 ( .A(n2029), .B(n1901), .CI(n1084), .CO(n1062), .S(n1063) );
  FA_X1 U752 ( .A(n2061), .B(n1869), .CI(n1837), .CO(n1064), .S(n1065) );
  FA_X1 U753 ( .A(n1773), .B(n1742), .CI(n1805), .CO(n1066), .S(n1067) );
  FA_X1 U754 ( .A(n1088), .B(n1073), .CI(n1071), .CO(n1068), .S(n1069) );
  FA_X1 U755 ( .A(n1075), .B(n1092), .CI(n1090), .CO(n1070), .S(n1071) );
  FA_X1 U756 ( .A(n1079), .B(n1094), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U757 ( .A(n1096), .B(n1098), .CI(n1081), .CO(n1074), .S(n1075) );
  FA_X1 U758 ( .A(n1085), .B(n1100), .CI(n1083), .CO(n1076), .S(n1077) );
  FA_X1 U759 ( .A(n1998), .B(n2062), .CI(n2030), .CO(n1078), .S(n1079) );
  FA_X1 U760 ( .A(n1966), .B(n1870), .CI(n1934), .CO(n1080), .S(n1081) );
  FA_X1 U761 ( .A(n1102), .B(n1838), .CI(n1902), .CO(n1082), .S(n1083) );
  FA_X1 U762 ( .A(n1774), .B(n1743), .CI(n1806), .CO(n1084), .S(n1085) );
  FA_X1 U763 ( .A(n1106), .B(n1091), .CI(n1089), .CO(n1086), .S(n1087) );
  FA_X1 U764 ( .A(n1108), .B(n1110), .CI(n1093), .CO(n1088), .S(n1089) );
  FA_X1 U765 ( .A(n1097), .B(n1099), .CI(n1095), .CO(n1090), .S(n1091) );
  FA_X1 U766 ( .A(n1114), .B(n1116), .CI(n1112), .CO(n1092), .S(n1093) );
  FA_X1 U767 ( .A(n1118), .B(n1999), .CI(n1101), .CO(n1094), .S(n1095) );
  FA_X1 U768 ( .A(n2063), .B(n1935), .CI(n2031), .CO(n1096), .S(n1097) );
  FA_X1 U769 ( .A(n1903), .B(n1103), .CI(n1967), .CO(n1098), .S(n1099) );
  FA_X1 U770 ( .A(n1871), .B(n1807), .CI(n1839), .CO(n1100), .S(n1101) );
  FA_X1 U771 ( .A(n1775), .B(n1744), .CI(n1120), .CO(n1102), .S(n1103) );
  FA_X1 U772 ( .A(n1124), .B(n1109), .CI(n1107), .CO(n1104), .S(n1105) );
  FA_X1 U773 ( .A(n1126), .B(n1128), .CI(n1111), .CO(n1106), .S(n1107) );
  FA_X1 U774 ( .A(n1115), .B(n1117), .CI(n1113), .CO(n1108), .S(n1109) );
  FA_X1 U775 ( .A(n1132), .B(n1119), .CI(n1130), .CO(n1110), .S(n1111) );
  FA_X1 U776 ( .A(n2064), .B(n2000), .CI(n1134), .CO(n1112), .S(n1113) );
  FA_X1 U777 ( .A(n2032), .B(n1936), .CI(n1136), .CO(n1114), .S(n1115) );
  FA_X1 U778 ( .A(n1872), .B(n1904), .CI(n1968), .CO(n1116), .S(n1117) );
  FA_X1 U779 ( .A(n1808), .B(n1121), .CI(n1840), .CO(n1118), .S(n1119) );
  HA_X1 U780 ( .A(n1776), .B(n1138), .CO(n1120), .S(n1121) );
  FA_X1 U781 ( .A(n1142), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U782 ( .A(n1129), .B(n1146), .CI(n1144), .CO(n1124), .S(n1125) );
  FA_X1 U783 ( .A(n1133), .B(n1148), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U784 ( .A(n1135), .B(n1137), .CI(n1150), .CO(n1128), .S(n1129) );
  FA_X1 U785 ( .A(n2033), .B(n2065), .CI(n1152), .CO(n1130), .S(n1131) );
  FA_X1 U786 ( .A(n2001), .B(n1905), .CI(n1969), .CO(n1132), .S(n1133) );
  FA_X1 U787 ( .A(n1154), .B(n1873), .CI(n1937), .CO(n1134), .S(n1135) );
  FA_X1 U788 ( .A(n1139), .B(n1809), .CI(n1841), .CO(n1136), .S(n1137) );
  HA_X1 U789 ( .A(n1156), .B(n1777), .CO(n1138), .S(n1139) );
  FA_X1 U790 ( .A(n1160), .B(n1145), .CI(n1143), .CO(n1140), .S(n1141) );
  FA_X1 U791 ( .A(n1147), .B(n1149), .CI(n1162), .CO(n1142), .S(n1143) );
  FA_X1 U792 ( .A(n1164), .B(n1166), .CI(n1151), .CO(n1144), .S(n1145) );
  FA_X1 U793 ( .A(n1153), .B(n2002), .CI(n1168), .CO(n1146), .S(n1147) );
  FA_X1 U794 ( .A(n1170), .B(n2034), .CI(n2066), .CO(n1148), .S(n1149) );
  FA_X1 U795 ( .A(n1938), .B(n1155), .CI(n1970), .CO(n1150), .S(n1151) );
  FA_X1 U796 ( .A(n1874), .B(n1842), .CI(n1906), .CO(n1152), .S(n1153) );
  FA_X1 U797 ( .A(n1810), .B(n1157), .CI(n1172), .CO(n1154), .S(n1155) );
  HA_X1 U798 ( .A(n289), .B(n1778), .CO(n1156), .S(n1157) );
  FA_X1 U799 ( .A(n1176), .B(n1163), .CI(n1161), .CO(n1158), .S(n1159) );
  FA_X1 U800 ( .A(n1165), .B(n1167), .CI(n1178), .CO(n1160), .S(n1161) );
  FA_X1 U801 ( .A(n1169), .B(n1182), .CI(n1180), .CO(n1162), .S(n1163) );
  FA_X1 U802 ( .A(n1184), .B(n2003), .CI(n1171), .CO(n1164), .S(n1165) );
  FA_X1 U803 ( .A(n2067), .B(n2035), .CI(n1186), .CO(n1166), .S(n1167) );
  FA_X1 U804 ( .A(n1907), .B(n1939), .CI(n1971), .CO(n1168), .S(n1169) );
  FA_X1 U805 ( .A(n1843), .B(n1173), .CI(n1875), .CO(n1170), .S(n1171) );
  HA_X1 U806 ( .A(n1811), .B(n1188), .CO(n1172), .S(n1173) );
  FA_X1 U807 ( .A(n1192), .B(n1179), .CI(n1177), .CO(n1174), .S(n1175) );
  FA_X1 U808 ( .A(n1181), .B(n1183), .CI(n1194), .CO(n1176), .S(n1177) );
  FA_X1 U809 ( .A(n1198), .B(n1185), .CI(n1196), .CO(n1178), .S(n1179) );
  FA_X1 U810 ( .A(n1200), .B(n2068), .CI(n1187), .CO(n1180), .S(n1181) );
  FA_X1 U811 ( .A(n2004), .B(n1940), .CI(n2036), .CO(n1182), .S(n1183) );
  FA_X1 U812 ( .A(n1202), .B(n1908), .CI(n1972), .CO(n1184), .S(n1185) );
  FA_X1 U813 ( .A(n1189), .B(n1844), .CI(n1876), .CO(n1186), .S(n1187) );
  HA_X1 U814 ( .A(n1204), .B(n1812), .CO(n1188), .S(n1189) );
  FA_X1 U815 ( .A(n1208), .B(n1195), .CI(n1193), .CO(n1190), .S(n1191) );
  FA_X1 U816 ( .A(n1197), .B(n1199), .CI(n1210), .CO(n1192), .S(n1193) );
  FA_X1 U817 ( .A(n1214), .B(n1201), .CI(n1212), .CO(n1194), .S(n1195) );
  FA_X1 U818 ( .A(n2037), .B(n2069), .CI(n1216), .CO(n1196), .S(n1197) );
  FA_X1 U819 ( .A(n1973), .B(n1203), .CI(n2005), .CO(n1198), .S(n1199) );
  FA_X1 U820 ( .A(n1941), .B(n1877), .CI(n1909), .CO(n1200), .S(n1201) );
  FA_X1 U821 ( .A(n1845), .B(n1205), .CI(n1218), .CO(n1202), .S(n1203) );
  HA_X1 U822 ( .A(n286), .B(n1813), .CO(n1204), .S(n1205) );
  FA_X1 U823 ( .A(n1222), .B(n1211), .CI(n1209), .CO(n1206), .S(n1207) );
  FA_X1 U824 ( .A(n1213), .B(n1215), .CI(n1224), .CO(n1208), .S(n1209) );
  FA_X1 U825 ( .A(n1217), .B(n1228), .CI(n1226), .CO(n1210), .S(n1211) );
  FA_X1 U826 ( .A(n2038), .B(n2070), .CI(n1230), .CO(n1212), .S(n1213) );
  FA_X1 U827 ( .A(n1942), .B(n1974), .CI(n2006), .CO(n1214), .S(n1215) );
  FA_X1 U828 ( .A(n1878), .B(n1219), .CI(n1910), .CO(n1216), .S(n1217) );
  HA_X1 U829 ( .A(n1846), .B(n1232), .CO(n1218), .S(n1219) );
  FA_X1 U830 ( .A(n1236), .B(n1225), .CI(n1223), .CO(n1220), .S(n1221) );
  FA_X1 U831 ( .A(n1227), .B(n1240), .CI(n1238), .CO(n1222), .S(n1223) );
  FA_X1 U832 ( .A(n1231), .B(n1242), .CI(n1229), .CO(n1224), .S(n1225) );
  FA_X1 U833 ( .A(n2071), .B(n1975), .CI(n2039), .CO(n1226), .S(n1227) );
  FA_X1 U834 ( .A(n1244), .B(n1943), .CI(n2007), .CO(n1228), .S(n1229) );
  FA_X1 U835 ( .A(n1233), .B(n1879), .CI(n1911), .CO(n1230), .S(n1231) );
  HA_X1 U836 ( .A(n1246), .B(n1847), .CO(n1232), .S(n1233) );
  FA_X1 U837 ( .A(n1250), .B(n1239), .CI(n1237), .CO(n1234), .S(n1235) );
  FA_X1 U838 ( .A(n1252), .B(n1254), .CI(n1241), .CO(n1236), .S(n1237) );
  FA_X1 U839 ( .A(n1256), .B(n2040), .CI(n1243), .CO(n1238), .S(n1239) );
  FA_X1 U840 ( .A(n2008), .B(n1245), .CI(n2072), .CO(n1240), .S(n1241) );
  FA_X1 U841 ( .A(n1944), .B(n1912), .CI(n1976), .CO(n1242), .S(n1243) );
  FA_X1 U842 ( .A(n1880), .B(n1247), .CI(n1258), .CO(n1244), .S(n1245) );
  HA_X1 U843 ( .A(n283), .B(n1848), .CO(n1246), .S(n1247) );
  FA_X1 U844 ( .A(n1262), .B(n1253), .CI(n1251), .CO(n1248), .S(n1249) );
  FA_X1 U845 ( .A(n1264), .B(n1257), .CI(n1255), .CO(n1250), .S(n1251) );
  FA_X1 U846 ( .A(n1268), .B(n2041), .CI(n1266), .CO(n1252), .S(n1253) );
  FA_X1 U847 ( .A(n1977), .B(n2009), .CI(n2073), .CO(n1254), .S(n1255) );
  FA_X1 U848 ( .A(n1913), .B(n1259), .CI(n1945), .CO(n1256), .S(n1257) );
  HA_X1 U849 ( .A(n1881), .B(n1270), .CO(n1258), .S(n1259) );
  FA_X1 U850 ( .A(n1274), .B(n1265), .CI(n1263), .CO(n1260), .S(n1261) );
  FA_X1 U851 ( .A(n1267), .B(n1269), .CI(n1276), .CO(n1262), .S(n1263) );
  FA_X1 U852 ( .A(n2074), .B(n2010), .CI(n1278), .CO(n1264), .S(n1265) );
  FA_X1 U853 ( .A(n1280), .B(n1978), .CI(n2042), .CO(n1266), .S(n1267) );
  FA_X1 U854 ( .A(n1271), .B(n1914), .CI(n1946), .CO(n1268), .S(n1269) );
  HA_X1 U855 ( .A(n1282), .B(n1882), .CO(n1270), .S(n1271) );
  FA_X1 U856 ( .A(n1277), .B(n1286), .CI(n1275), .CO(n1272), .S(n1273) );
  FA_X1 U857 ( .A(n1279), .B(n1290), .CI(n1288), .CO(n1274), .S(n1275) );
  FA_X1 U858 ( .A(n2043), .B(n1281), .CI(n2075), .CO(n1276), .S(n1277) );
  FA_X1 U859 ( .A(n2011), .B(n1947), .CI(n1979), .CO(n1278), .S(n1279) );
  FA_X1 U860 ( .A(n1915), .B(n1283), .CI(n1292), .CO(n1280), .S(n1281) );
  HA_X1 U861 ( .A(n280), .B(n1883), .CO(n1282), .S(n1283) );
  FA_X1 U862 ( .A(n1296), .B(n1289), .CI(n1287), .CO(n1284), .S(n1285) );
  FA_X1 U863 ( .A(n1298), .B(n1300), .CI(n1291), .CO(n1286), .S(n1287) );
  FA_X1 U864 ( .A(n2012), .B(n2044), .CI(n2076), .CO(n1288), .S(n1289) );
  FA_X1 U865 ( .A(n1948), .B(n1293), .CI(n1980), .CO(n1290), .S(n1291) );
  HA_X1 U866 ( .A(n1916), .B(n1302), .CO(n1292), .S(n1293) );
  FA_X1 U867 ( .A(n1306), .B(n1299), .CI(n1297), .CO(n1294), .S(n1295) );
  FA_X1 U868 ( .A(n1308), .B(n2045), .CI(n1301), .CO(n1296), .S(n1297) );
  FA_X1 U869 ( .A(n1310), .B(n2013), .CI(n2077), .CO(n1298), .S(n1299) );
  FA_X1 U870 ( .A(n1303), .B(n1949), .CI(n1981), .CO(n1300), .S(n1301) );
  HA_X1 U871 ( .A(n1312), .B(n1917), .CO(n1302), .S(n1303) );
  FA_X1 U872 ( .A(n1316), .B(n1309), .CI(n1307), .CO(n1304), .S(n1305) );
  FA_X1 U873 ( .A(n2078), .B(n1311), .CI(n1318), .CO(n1306), .S(n1307) );
  FA_X1 U874 ( .A(n2046), .B(n1982), .CI(n2014), .CO(n1308), .S(n1309) );
  FA_X1 U875 ( .A(n1950), .B(n1313), .CI(n1320), .CO(n1310), .S(n1311) );
  HA_X1 U876 ( .A(n277), .B(n1918), .CO(n1312), .S(n1313) );
  FA_X1 U877 ( .A(n1324), .B(n1319), .CI(n1317), .CO(n1314), .S(n1315) );
  FA_X1 U878 ( .A(n2047), .B(n2079), .CI(n1326), .CO(n1316), .S(n1317) );
  FA_X1 U879 ( .A(n1983), .B(n1321), .CI(n2015), .CO(n1318), .S(n1319) );
  HA_X1 U880 ( .A(n1951), .B(n1328), .CO(n1320), .S(n1321) );
  FA_X1 U881 ( .A(n1327), .B(n1332), .CI(n1325), .CO(n1322), .S(n1323) );
  FA_X1 U882 ( .A(n1334), .B(n2048), .CI(n2080), .CO(n1324), .S(n1325) );
  FA_X1 U883 ( .A(n1329), .B(n1984), .CI(n2016), .CO(n1326), .S(n1327) );
  HA_X1 U884 ( .A(n1336), .B(n1952), .CO(n1328), .S(n1329) );
  FA_X1 U885 ( .A(n1340), .B(n1335), .CI(n1333), .CO(n1330), .S(n1331) );
  FA_X1 U886 ( .A(n2081), .B(n2017), .CI(n2049), .CO(n1332), .S(n1333) );
  FA_X1 U887 ( .A(n1985), .B(n1337), .CI(n1342), .CO(n1334), .S(n1335) );
  HA_X1 U888 ( .A(n274), .B(n1953), .CO(n1336), .S(n1337) );
  FA_X1 U889 ( .A(n1346), .B(n2082), .CI(n1341), .CO(n1338), .S(n1339) );
  FA_X1 U890 ( .A(n2018), .B(n1343), .CI(n2050), .CO(n1340), .S(n1341) );
  HA_X1 U891 ( .A(n1986), .B(n1348), .CO(n1342), .S(n1343) );
  FA_X1 U892 ( .A(n1352), .B(n2083), .CI(n1347), .CO(n1344), .S(n1345) );
  FA_X1 U893 ( .A(n1349), .B(n2019), .CI(n2051), .CO(n1346), .S(n1347) );
  HA_X1 U894 ( .A(n1354), .B(n1987), .CO(n1348), .S(n1349) );
  FA_X1 U895 ( .A(n2084), .B(n2052), .CI(n1353), .CO(n1350), .S(n1351) );
  FA_X1 U896 ( .A(n2020), .B(n1355), .CI(n1358), .CO(n1352), .S(n1353) );
  HA_X1 U897 ( .A(n271), .B(n1988), .CO(n1354), .S(n1355) );
  FA_X1 U898 ( .A(n2053), .B(n1359), .CI(n2085), .CO(n1356), .S(n1357) );
  HA_X1 U899 ( .A(n2021), .B(n1362), .CO(n1358), .S(n1359) );
  FA_X1 U900 ( .A(n1363), .B(n2054), .CI(n2086), .CO(n1360), .S(n1361) );
  HA_X1 U901 ( .A(n1366), .B(n2022), .CO(n1362), .S(n1363) );
  FA_X1 U902 ( .A(n2055), .B(n1367), .CI(n1368), .CO(n1364), .S(n1365) );
  HA_X1 U903 ( .A(n268), .B(n2023), .CO(n1366), .S(n1367) );
  HA_X1 U904 ( .A(n2056), .B(n1370), .CO(n1368), .S(n1369) );
  HA_X1 U905 ( .A(n1372), .B(n2057), .CO(n1370), .S(n1371) );
  HA_X1 U906 ( .A(n265), .B(n2058), .CO(n1372), .S(n1373) );
  OAI21_X4 U907 ( .B1(n2808), .B2(n366), .A(n2094), .ZN(n1720) );
  NAND2_X4 U908 ( .A1(n388), .A2(n484), .ZN(n2094) );
  OAI21_X4 U909 ( .B1(n2809), .B2(n366), .A(n2095), .ZN(n717) );
  AOI21_X4 U910 ( .B1(n388), .B2(n481), .A(n1374), .ZN(n2095) );
  AND2_X4 U911 ( .A1(n333), .A2(n484), .ZN(n1374) );
  OAI21_X4 U912 ( .B1(n2810), .B2(n366), .A(n2096), .ZN(n1721) );
  AOI222_X2 U913 ( .A1(n3131), .A2(n484), .B1(n333), .B2(n481), .C1(n388), 
        .C2(n478), .ZN(n2096) );
  OAI21_X4 U914 ( .B1(n2811), .B2(n366), .A(n2097), .ZN(n1722) );
  AOI222_X2 U915 ( .A1(n3130), .A2(n481), .B1(n333), .B2(n478), .C1(n388), 
        .C2(n475), .ZN(n2097) );
  OAI21_X4 U916 ( .B1(n2812), .B2(n366), .A(n2098), .ZN(n723) );
  AOI222_X2 U917 ( .A1(n3131), .A2(n478), .B1(n333), .B2(n475), .C1(n388), 
        .C2(n472), .ZN(n2098) );
  OAI21_X4 U918 ( .B1(n2813), .B2(n366), .A(n2099), .ZN(n1723) );
  AOI222_X2 U919 ( .A1(n3130), .A2(n475), .B1(n333), .B2(n472), .C1(n388), 
        .C2(n469), .ZN(n2099) );
  OAI21_X4 U920 ( .B1(n2814), .B2(n366), .A(n2100), .ZN(n1724) );
  AOI222_X2 U921 ( .A1(n3131), .A2(n472), .B1(n333), .B2(n469), .C1(n388), 
        .C2(n466), .ZN(n2100) );
  OAI21_X4 U922 ( .B1(n2815), .B2(n366), .A(n2101), .ZN(n736) );
  AOI222_X2 U923 ( .A1(n3130), .A2(n469), .B1(n333), .B2(n466), .C1(n388), 
        .C2(n463), .ZN(n2101) );
  OAI21_X4 U924 ( .B1(n2816), .B2(n366), .A(n2102), .ZN(n1725) );
  AOI222_X2 U925 ( .A1(n3131), .A2(n466), .B1(n333), .B2(n463), .C1(n388), 
        .C2(n460), .ZN(n2102) );
  OAI21_X4 U926 ( .B1(n2817), .B2(n366), .A(n2103), .ZN(n1726) );
  AOI222_X2 U927 ( .A1(n3130), .A2(n463), .B1(n333), .B2(n460), .C1(n388), 
        .C2(n457), .ZN(n2103) );
  OAI21_X4 U928 ( .B1(n2818), .B2(n366), .A(n2104), .ZN(n755) );
  AOI222_X2 U929 ( .A1(n3131), .A2(n460), .B1(n333), .B2(n457), .C1(n388), 
        .C2(n454), .ZN(n2104) );
  OAI21_X4 U930 ( .B1(n2819), .B2(n366), .A(n2105), .ZN(n1727) );
  AOI222_X2 U931 ( .A1(n3130), .A2(n457), .B1(n333), .B2(n454), .C1(n388), 
        .C2(n451), .ZN(n2105) );
  OAI21_X4 U932 ( .B1(n2820), .B2(n366), .A(n2106), .ZN(n1728) );
  AOI222_X2 U933 ( .A1(n3131), .A2(n454), .B1(n333), .B2(n451), .C1(n388), 
        .C2(n448), .ZN(n2106) );
  OAI21_X4 U934 ( .B1(n2821), .B2(n366), .A(n2107), .ZN(n780) );
  AOI222_X2 U935 ( .A1(n3130), .A2(n451), .B1(n333), .B2(n448), .C1(n388), 
        .C2(n445), .ZN(n2107) );
  OAI21_X4 U936 ( .B1(n2822), .B2(n366), .A(n2108), .ZN(n1729) );
  AOI222_X2 U937 ( .A1(n3131), .A2(n448), .B1(n333), .B2(n445), .C1(n388), 
        .C2(n442), .ZN(n2108) );
  OAI21_X4 U938 ( .B1(n2823), .B2(n366), .A(n2109), .ZN(n1730) );
  AOI222_X2 U939 ( .A1(n3130), .A2(n445), .B1(n333), .B2(n442), .C1(n388), 
        .C2(n439), .ZN(n2109) );
  OAI21_X4 U940 ( .B1(n2824), .B2(n366), .A(n2110), .ZN(n811) );
  AOI222_X2 U941 ( .A1(n3131), .A2(n442), .B1(n333), .B2(n439), .C1(n388), 
        .C2(n436), .ZN(n2110) );
  OAI21_X4 U942 ( .B1(n2825), .B2(n366), .A(n2111), .ZN(n1731) );
  AOI222_X2 U943 ( .A1(n3130), .A2(n439), .B1(n333), .B2(n436), .C1(n388), 
        .C2(n433), .ZN(n2111) );
  OAI21_X4 U944 ( .B1(n2826), .B2(n366), .A(n2112), .ZN(n1732) );
  AOI222_X2 U945 ( .A1(n3131), .A2(n436), .B1(n333), .B2(n433), .C1(n388), 
        .C2(n430), .ZN(n2112) );
  OAI21_X4 U946 ( .B1(n2827), .B2(n366), .A(n2113), .ZN(n848) );
  AOI222_X2 U947 ( .A1(n3130), .A2(n433), .B1(n333), .B2(n430), .C1(n388), 
        .C2(n427), .ZN(n2113) );
  OAI21_X4 U948 ( .B1(n2828), .B2(n366), .A(n2114), .ZN(n1733) );
  AOI222_X2 U949 ( .A1(n3131), .A2(n430), .B1(n333), .B2(n427), .C1(n388), 
        .C2(n424), .ZN(n2114) );
  OAI21_X4 U950 ( .B1(n2829), .B2(n366), .A(n2115), .ZN(n891) );
  AOI222_X2 U951 ( .A1(n3130), .A2(n427), .B1(n333), .B2(n424), .C1(n388), 
        .C2(n421), .ZN(n2115) );
  OAI21_X4 U952 ( .B1(n2830), .B2(n366), .A(n2116), .ZN(n1734) );
  AOI222_X2 U953 ( .A1(n3131), .A2(n424), .B1(n333), .B2(n421), .C1(n388), 
        .C2(n418), .ZN(n2116) );
  OAI21_X4 U954 ( .B1(n2831), .B2(n366), .A(n2117), .ZN(n1735) );
  AOI222_X2 U955 ( .A1(n3131), .A2(n421), .B1(n333), .B2(n418), .C1(n388), 
        .C2(n415), .ZN(n2117) );
  OAI21_X4 U956 ( .B1(n2832), .B2(n366), .A(n2118), .ZN(n1736) );
  AOI222_X2 U957 ( .A1(n3130), .A2(n418), .B1(n333), .B2(n415), .C1(n388), 
        .C2(n412), .ZN(n2118) );
  OAI21_X4 U958 ( .B1(n2833), .B2(n366), .A(n2119), .ZN(n941) );
  AOI222_X2 U959 ( .A1(n3130), .A2(n415), .B1(n333), .B2(n412), .C1(n388), 
        .C2(n409), .ZN(n2119) );
  AOI222_X2 U961 ( .A1(n3131), .A2(n412), .B1(n333), .B2(n409), .C1(n388), 
        .C2(n406), .ZN(n2120) );
  OAI21_X4 U962 ( .B1(n2835), .B2(n366), .A(n2121), .ZN(n1738) );
  AOI222_X2 U963 ( .A1(n3130), .A2(n409), .B1(n333), .B2(n406), .C1(n388), 
        .C2(n403), .ZN(n2121) );
  OAI21_X4 U964 ( .B1(n2836), .B2(n366), .A(n2122), .ZN(n1739) );
  AOI222_X2 U965 ( .A1(n3131), .A2(n406), .B1(n333), .B2(n403), .C1(n388), 
        .C2(n400), .ZN(n2122) );
  OAI21_X4 U966 ( .B1(n2837), .B2(n366), .A(n2123), .ZN(n1740) );
  AOI222_X2 U967 ( .A1(n3130), .A2(n403), .B1(n333), .B2(n400), .C1(n388), 
        .C2(n397), .ZN(n2123) );
  OAI21_X4 U968 ( .B1(n2838), .B2(n366), .A(n2124), .ZN(n1741) );
  AOI222_X2 U969 ( .A1(n3131), .A2(n400), .B1(n333), .B2(n397), .C1(n388), 
        .C2(n393), .ZN(n2124) );
  OAI21_X4 U970 ( .B1(n2839), .B2(n366), .A(n2125), .ZN(n1742) );
  AOI222_X2 U971 ( .A1(n3131), .A2(n397), .B1(n333), .B2(n393), .C1(n388), 
        .C2(n390), .ZN(n2125) );
  OAI21_X4 U972 ( .B1(n2840), .B2(n366), .A(n2126), .ZN(n1743) );
  OAI21_X4 U974 ( .B1(n2841), .B2(n366), .A(n2127), .ZN(n1744) );
  AND2_X4 U976 ( .A1(n3130), .A2(n390), .ZN(n1376) );
  XOR2_X2 U978 ( .A(n2128), .B(n289), .Z(n1746) );
  OAI21_X4 U979 ( .B1(n2808), .B2(n363), .A(n2162), .ZN(n2128) );
  NAND2_X4 U980 ( .A1(n386), .A2(n484), .ZN(n2162) );
  XOR2_X2 U981 ( .A(n2129), .B(n289), .Z(n1747) );
  OAI21_X4 U982 ( .B1(n2809), .B2(n363), .A(n2163), .ZN(n2129) );
  AOI21_X4 U983 ( .B1(n386), .B2(n481), .A(n1377), .ZN(n2163) );
  AND2_X4 U984 ( .A1(n331), .A2(n484), .ZN(n1377) );
  XOR2_X2 U985 ( .A(n2130), .B(n289), .Z(n1748) );
  OAI21_X4 U986 ( .B1(n2810), .B2(n363), .A(n2164), .ZN(n2130) );
  AOI222_X2 U987 ( .A1(n3128), .A2(n484), .B1(n331), .B2(n481), .C1(n386), 
        .C2(n478), .ZN(n2164) );
  XOR2_X2 U988 ( .A(n2131), .B(n289), .Z(n1749) );
  OAI21_X4 U989 ( .B1(n2811), .B2(n363), .A(n2165), .ZN(n2131) );
  AOI222_X2 U990 ( .A1(n3127), .A2(n481), .B1(n331), .B2(n478), .C1(n386), 
        .C2(n475), .ZN(n2165) );
  XOR2_X2 U991 ( .A(n2132), .B(n289), .Z(n1750) );
  OAI21_X4 U992 ( .B1(n2812), .B2(n363), .A(n2166), .ZN(n2132) );
  AOI222_X2 U993 ( .A1(n3128), .A2(n478), .B1(n331), .B2(n475), .C1(n386), 
        .C2(n472), .ZN(n2166) );
  XOR2_X2 U994 ( .A(n2133), .B(n289), .Z(n1751) );
  OAI21_X4 U995 ( .B1(n2813), .B2(n363), .A(n2167), .ZN(n2133) );
  AOI222_X2 U996 ( .A1(n3127), .A2(n475), .B1(n331), .B2(n472), .C1(n386), 
        .C2(n469), .ZN(n2167) );
  XOR2_X2 U997 ( .A(n2134), .B(n289), .Z(n1752) );
  OAI21_X4 U998 ( .B1(n2814), .B2(n363), .A(n2168), .ZN(n2134) );
  AOI222_X2 U999 ( .A1(n3128), .A2(n472), .B1(n331), .B2(n469), .C1(n386), 
        .C2(n466), .ZN(n2168) );
  XOR2_X2 U1000 ( .A(n2135), .B(n289), .Z(n1753) );
  OAI21_X4 U1001 ( .B1(n2815), .B2(n363), .A(n2169), .ZN(n2135) );
  AOI222_X2 U1002 ( .A1(n3127), .A2(n469), .B1(n331), .B2(n466), .C1(n386), 
        .C2(n463), .ZN(n2169) );
  XOR2_X2 U1003 ( .A(n2136), .B(n289), .Z(n1754) );
  OAI21_X4 U1004 ( .B1(n2816), .B2(n363), .A(n2170), .ZN(n2136) );
  AOI222_X2 U1005 ( .A1(n3128), .A2(n466), .B1(n331), .B2(n463), .C1(n386), 
        .C2(n460), .ZN(n2170) );
  XOR2_X2 U1006 ( .A(n2137), .B(n289), .Z(n1755) );
  OAI21_X4 U1007 ( .B1(n2817), .B2(n363), .A(n2171), .ZN(n2137) );
  AOI222_X2 U1008 ( .A1(n3127), .A2(n463), .B1(n331), .B2(n460), .C1(n386), 
        .C2(n457), .ZN(n2171) );
  XOR2_X2 U1009 ( .A(n2138), .B(n289), .Z(n1756) );
  OAI21_X4 U1010 ( .B1(n2818), .B2(n363), .A(n2172), .ZN(n2138) );
  AOI222_X2 U1011 ( .A1(n3128), .A2(n460), .B1(n331), .B2(n457), .C1(n386), 
        .C2(n454), .ZN(n2172) );
  XOR2_X2 U1012 ( .A(n2139), .B(n289), .Z(n1757) );
  OAI21_X4 U1013 ( .B1(n2819), .B2(n363), .A(n2173), .ZN(n2139) );
  AOI222_X2 U1014 ( .A1(n3127), .A2(n457), .B1(n331), .B2(n454), .C1(n386), 
        .C2(n451), .ZN(n2173) );
  XOR2_X2 U1015 ( .A(n2140), .B(n289), .Z(n1758) );
  OAI21_X4 U1016 ( .B1(n2820), .B2(n363), .A(n2174), .ZN(n2140) );
  AOI222_X2 U1017 ( .A1(n3127), .A2(n454), .B1(n331), .B2(n451), .C1(n386), 
        .C2(n448), .ZN(n2174) );
  XOR2_X2 U1018 ( .A(n2141), .B(n289), .Z(n1759) );
  OAI21_X4 U1019 ( .B1(n2821), .B2(n363), .A(n2175), .ZN(n2141) );
  AOI222_X2 U1020 ( .A1(n3128), .A2(n451), .B1(n331), .B2(n448), .C1(n386), 
        .C2(n445), .ZN(n2175) );
  XOR2_X2 U1021 ( .A(n2142), .B(n289), .Z(n1760) );
  OAI21_X4 U1022 ( .B1(n2822), .B2(n363), .A(n2176), .ZN(n2142) );
  AOI222_X2 U1023 ( .A1(n3128), .A2(n448), .B1(n331), .B2(n445), .C1(n386), 
        .C2(n442), .ZN(n2176) );
  XOR2_X2 U1024 ( .A(n2143), .B(n289), .Z(n1761) );
  OAI21_X4 U1025 ( .B1(n2823), .B2(n363), .A(n2177), .ZN(n2143) );
  AOI222_X2 U1026 ( .A1(n3127), .A2(n445), .B1(n331), .B2(n442), .C1(n386), 
        .C2(n439), .ZN(n2177) );
  XOR2_X2 U1027 ( .A(n2144), .B(n289), .Z(n1762) );
  OAI21_X4 U1028 ( .B1(n2824), .B2(n363), .A(n2178), .ZN(n2144) );
  AOI222_X2 U1029 ( .A1(n3128), .A2(n442), .B1(n331), .B2(n439), .C1(n386), 
        .C2(n436), .ZN(n2178) );
  XOR2_X2 U1030 ( .A(n2145), .B(n289), .Z(n1763) );
  OAI21_X4 U1031 ( .B1(n2825), .B2(n363), .A(n2179), .ZN(n2145) );
  AOI222_X2 U1032 ( .A1(n3127), .A2(n439), .B1(n331), .B2(n436), .C1(n386), 
        .C2(n433), .ZN(n2179) );
  XOR2_X2 U1033 ( .A(n2146), .B(n289), .Z(n1764) );
  OAI21_X4 U1034 ( .B1(n2826), .B2(n363), .A(n2180), .ZN(n2146) );
  AOI222_X2 U1035 ( .A1(n3128), .A2(n436), .B1(n331), .B2(n433), .C1(n386), 
        .C2(n430), .ZN(n2180) );
  XOR2_X2 U1036 ( .A(n2147), .B(n289), .Z(n907) );
  OAI21_X4 U1037 ( .B1(n2827), .B2(n363), .A(n2181), .ZN(n2147) );
  AOI222_X2 U1038 ( .A1(n3127), .A2(n433), .B1(n331), .B2(n430), .C1(n386), 
        .C2(n427), .ZN(n2181) );
  XOR2_X2 U1039 ( .A(n2148), .B(n289), .Z(n1765) );
  OAI21_X4 U1040 ( .B1(n2828), .B2(n363), .A(n2182), .ZN(n2148) );
  AOI222_X2 U1041 ( .A1(n3128), .A2(n430), .B1(n331), .B2(n427), .C1(n386), 
        .C2(n424), .ZN(n2182) );
  XOR2_X2 U1042 ( .A(n2149), .B(n289), .Z(n1766) );
  OAI21_X4 U1043 ( .B1(n2829), .B2(n363), .A(n2183), .ZN(n2149) );
  AOI222_X2 U1044 ( .A1(n3127), .A2(n427), .B1(n331), .B2(n424), .C1(n386), 
        .C2(n421), .ZN(n2183) );
  XOR2_X2 U1045 ( .A(n2150), .B(n289), .Z(n1767) );
  OAI21_X4 U1046 ( .B1(n2830), .B2(n363), .A(n2184), .ZN(n2150) );
  AOI222_X2 U1047 ( .A1(n3128), .A2(n424), .B1(n331), .B2(n421), .C1(n386), 
        .C2(n418), .ZN(n2184) );
  XOR2_X2 U1048 ( .A(n2151), .B(n289), .Z(n1768) );
  OAI21_X4 U1049 ( .B1(n2831), .B2(n363), .A(n2185), .ZN(n2151) );
  AOI222_X2 U1050 ( .A1(n3127), .A2(n421), .B1(n331), .B2(n418), .C1(n386), 
        .C2(n415), .ZN(n2185) );
  XOR2_X2 U1051 ( .A(n2152), .B(n289), .Z(n1769) );
  OAI21_X4 U1052 ( .B1(n2832), .B2(n363), .A(n2186), .ZN(n2152) );
  AOI222_X2 U1053 ( .A1(n3128), .A2(n418), .B1(n331), .B2(n415), .C1(n386), 
        .C2(n412), .ZN(n2186) );
  XOR2_X2 U1054 ( .A(n2153), .B(n289), .Z(n1770) );
  OAI21_X4 U1055 ( .B1(n2833), .B2(n363), .A(n2187), .ZN(n2153) );
  AOI222_X2 U1056 ( .A1(n3127), .A2(n415), .B1(n331), .B2(n412), .C1(n386), 
        .C2(n409), .ZN(n2187) );
  XOR2_X2 U1057 ( .A(n2154), .B(n289), .Z(n1771) );
  AOI222_X2 U1059 ( .A1(n3128), .A2(n412), .B1(n331), .B2(n409), .C1(n386), 
        .C2(n406), .ZN(n2188) );
  XOR2_X2 U1060 ( .A(n2155), .B(n289), .Z(n1772) );
  OAI21_X4 U1061 ( .B1(n2835), .B2(n363), .A(n2189), .ZN(n2155) );
  AOI222_X2 U1062 ( .A1(n3127), .A2(n409), .B1(n331), .B2(n406), .C1(n386), 
        .C2(n403), .ZN(n2189) );
  XOR2_X2 U1063 ( .A(n2156), .B(n289), .Z(n1773) );
  OAI21_X4 U1064 ( .B1(n2836), .B2(n363), .A(n2190), .ZN(n2156) );
  AOI222_X2 U1065 ( .A1(n3128), .A2(n406), .B1(n331), .B2(n403), .C1(n386), 
        .C2(n400), .ZN(n2190) );
  XOR2_X2 U1066 ( .A(n2157), .B(n289), .Z(n1774) );
  OAI21_X4 U1067 ( .B1(n2837), .B2(n363), .A(n2191), .ZN(n2157) );
  AOI222_X2 U1068 ( .A1(n3127), .A2(n403), .B1(n331), .B2(n400), .C1(n386), 
        .C2(n397), .ZN(n2191) );
  XOR2_X2 U1069 ( .A(n2158), .B(n289), .Z(n1775) );
  OAI21_X4 U1070 ( .B1(n2838), .B2(n363), .A(n2192), .ZN(n2158) );
  AOI222_X2 U1071 ( .A1(n3128), .A2(n400), .B1(n331), .B2(n397), .C1(n386), 
        .C2(n393), .ZN(n2192) );
  XOR2_X2 U1072 ( .A(n2159), .B(n289), .Z(n1776) );
  OAI21_X4 U1073 ( .B1(n2839), .B2(n363), .A(n2193), .ZN(n2159) );
  AOI222_X2 U1074 ( .A1(n3127), .A2(n397), .B1(n331), .B2(n393), .C1(n386), 
        .C2(n390), .ZN(n2193) );
  XOR2_X2 U1075 ( .A(n2160), .B(n289), .Z(n1777) );
  OAI21_X4 U1076 ( .B1(n2840), .B2(n363), .A(n2194), .ZN(n2160) );
  XOR2_X2 U1078 ( .A(n2161), .B(n289), .Z(n1778) );
  OAI21_X4 U1079 ( .B1(n2841), .B2(n363), .A(n2195), .ZN(n2161) );
  AND2_X4 U1081 ( .A1(n3127), .A2(n390), .ZN(n1379) );
  XOR2_X2 U1083 ( .A(n2196), .B(n286), .Z(n1780) );
  OAI21_X4 U1084 ( .B1(n2808), .B2(n360), .A(n2230), .ZN(n2196) );
  NAND2_X4 U1085 ( .A1(n384), .A2(n484), .ZN(n2230) );
  XOR2_X2 U1086 ( .A(n2197), .B(n286), .Z(n1781) );
  OAI21_X4 U1087 ( .B1(n2809), .B2(n360), .A(n2231), .ZN(n2197) );
  AOI21_X4 U1088 ( .B1(n384), .B2(n481), .A(n1380), .ZN(n2231) );
  AND2_X4 U1089 ( .A1(n329), .A2(n484), .ZN(n1380) );
  XOR2_X2 U1090 ( .A(n2198), .B(n286), .Z(n1782) );
  OAI21_X4 U1091 ( .B1(n2810), .B2(n360), .A(n2232), .ZN(n2198) );
  AOI222_X2 U1092 ( .A1(n3141), .A2(n484), .B1(n329), .B2(n481), .C1(n384), 
        .C2(n478), .ZN(n2232) );
  XOR2_X2 U1093 ( .A(n2199), .B(n286), .Z(n1783) );
  OAI21_X4 U1094 ( .B1(n2811), .B2(n360), .A(n2233), .ZN(n2199) );
  AOI222_X2 U1095 ( .A1(n3141), .A2(n481), .B1(n329), .B2(n478), .C1(n384), 
        .C2(n475), .ZN(n2233) );
  XOR2_X2 U1096 ( .A(n2200), .B(n286), .Z(n1784) );
  OAI21_X4 U1097 ( .B1(n2812), .B2(n360), .A(n2234), .ZN(n2200) );
  AOI222_X2 U1098 ( .A1(n3141), .A2(n478), .B1(n329), .B2(n475), .C1(n384), 
        .C2(n472), .ZN(n2234) );
  XOR2_X2 U1099 ( .A(n2201), .B(n286), .Z(n1785) );
  OAI21_X4 U1100 ( .B1(n2813), .B2(n360), .A(n2235), .ZN(n2201) );
  AOI222_X2 U1101 ( .A1(n3141), .A2(n475), .B1(n329), .B2(n472), .C1(n384), 
        .C2(n469), .ZN(n2235) );
  XOR2_X2 U1102 ( .A(n2202), .B(n286), .Z(n1786) );
  OAI21_X4 U1103 ( .B1(n2814), .B2(n360), .A(n2236), .ZN(n2202) );
  AOI222_X2 U1104 ( .A1(n3141), .A2(n472), .B1(n329), .B2(n469), .C1(n384), 
        .C2(n466), .ZN(n2236) );
  XOR2_X2 U1105 ( .A(n2203), .B(n286), .Z(n1787) );
  OAI21_X4 U1106 ( .B1(n2815), .B2(n360), .A(n2237), .ZN(n2203) );
  AOI222_X2 U1107 ( .A1(n3141), .A2(n469), .B1(n329), .B2(n466), .C1(n384), 
        .C2(n463), .ZN(n2237) );
  XOR2_X2 U1108 ( .A(n2204), .B(n286), .Z(n1788) );
  OAI21_X4 U1109 ( .B1(n2816), .B2(n360), .A(n2238), .ZN(n2204) );
  AOI222_X2 U1110 ( .A1(n3141), .A2(n466), .B1(n329), .B2(n463), .C1(n384), 
        .C2(n460), .ZN(n2238) );
  XOR2_X2 U1111 ( .A(n2205), .B(n286), .Z(n1789) );
  OAI21_X4 U1112 ( .B1(n2817), .B2(n360), .A(n2239), .ZN(n2205) );
  AOI222_X2 U1113 ( .A1(n3141), .A2(n463), .B1(n329), .B2(n460), .C1(n384), 
        .C2(n457), .ZN(n2239) );
  XOR2_X2 U1114 ( .A(n2206), .B(n286), .Z(n1790) );
  OAI21_X4 U1115 ( .B1(n2818), .B2(n360), .A(n2240), .ZN(n2206) );
  AOI222_X2 U1116 ( .A1(n3141), .A2(n460), .B1(n329), .B2(n457), .C1(n384), 
        .C2(n454), .ZN(n2240) );
  XOR2_X2 U1117 ( .A(n2207), .B(n286), .Z(n1791) );
  OAI21_X4 U1118 ( .B1(n2819), .B2(n360), .A(n2241), .ZN(n2207) );
  AOI222_X2 U1119 ( .A1(n3141), .A2(n457), .B1(n329), .B2(n454), .C1(n384), 
        .C2(n451), .ZN(n2241) );
  XOR2_X2 U1120 ( .A(n2208), .B(n286), .Z(n1792) );
  OAI21_X4 U1121 ( .B1(n2820), .B2(n360), .A(n2242), .ZN(n2208) );
  AOI222_X2 U1122 ( .A1(n3141), .A2(n454), .B1(n329), .B2(n451), .C1(n384), 
        .C2(n448), .ZN(n2242) );
  XOR2_X2 U1123 ( .A(n2209), .B(n286), .Z(n1793) );
  OAI21_X4 U1124 ( .B1(n2821), .B2(n360), .A(n2243), .ZN(n2209) );
  AOI222_X2 U1125 ( .A1(n3141), .A2(n451), .B1(n329), .B2(n448), .C1(n384), 
        .C2(n445), .ZN(n2243) );
  XOR2_X2 U1126 ( .A(n2210), .B(n286), .Z(n1794) );
  OAI21_X4 U1127 ( .B1(n2822), .B2(n360), .A(n2244), .ZN(n2210) );
  AOI222_X2 U1128 ( .A1(n3141), .A2(n448), .B1(n329), .B2(n445), .C1(n384), 
        .C2(n442), .ZN(n2244) );
  XOR2_X2 U1129 ( .A(n2211), .B(n286), .Z(n1795) );
  OAI21_X4 U1130 ( .B1(n2823), .B2(n360), .A(n2245), .ZN(n2211) );
  AOI222_X2 U1131 ( .A1(n3141), .A2(n445), .B1(n329), .B2(n442), .C1(n384), 
        .C2(n439), .ZN(n2245) );
  XOR2_X2 U1132 ( .A(n2212), .B(n286), .Z(n1796) );
  OAI21_X4 U1133 ( .B1(n2824), .B2(n360), .A(n2246), .ZN(n2212) );
  AOI222_X2 U1134 ( .A1(n3141), .A2(n442), .B1(n329), .B2(n439), .C1(n384), 
        .C2(n436), .ZN(n2246) );
  XOR2_X2 U1135 ( .A(n2213), .B(n286), .Z(n1797) );
  OAI21_X4 U1136 ( .B1(n2825), .B2(n360), .A(n2247), .ZN(n2213) );
  AOI222_X2 U1137 ( .A1(n3141), .A2(n439), .B1(n329), .B2(n436), .C1(n384), 
        .C2(n433), .ZN(n2247) );
  XOR2_X2 U1138 ( .A(n2214), .B(n286), .Z(n1798) );
  OAI21_X4 U1139 ( .B1(n2826), .B2(n360), .A(n2248), .ZN(n2214) );
  AOI222_X2 U1140 ( .A1(n3141), .A2(n436), .B1(n329), .B2(n433), .C1(n384), 
        .C2(n430), .ZN(n2248) );
  XOR2_X2 U1141 ( .A(n2215), .B(n286), .Z(n1799) );
  OAI21_X4 U1142 ( .B1(n2827), .B2(n360), .A(n2249), .ZN(n2215) );
  AOI222_X2 U1143 ( .A1(n3141), .A2(n433), .B1(n329), .B2(n430), .C1(n384), 
        .C2(n427), .ZN(n2249) );
  XOR2_X2 U1144 ( .A(n2216), .B(n286), .Z(n1800) );
  OAI21_X4 U1145 ( .B1(n2828), .B2(n360), .A(n2250), .ZN(n2216) );
  AOI222_X2 U1146 ( .A1(n3141), .A2(n430), .B1(n329), .B2(n427), .C1(n384), 
        .C2(n424), .ZN(n2250) );
  XOR2_X2 U1147 ( .A(n2217), .B(n286), .Z(n1801) );
  OAI21_X4 U1148 ( .B1(n2829), .B2(n360), .A(n2251), .ZN(n2217) );
  AOI222_X2 U1149 ( .A1(n3141), .A2(n427), .B1(n329), .B2(n424), .C1(n384), 
        .C2(n421), .ZN(n2251) );
  XOR2_X2 U1150 ( .A(n2218), .B(n286), .Z(n1802) );
  OAI21_X4 U1151 ( .B1(n2830), .B2(n360), .A(n2252), .ZN(n2218) );
  AOI222_X2 U1152 ( .A1(n3141), .A2(n424), .B1(n329), .B2(n421), .C1(n384), 
        .C2(n418), .ZN(n2252) );
  XOR2_X2 U1153 ( .A(n2219), .B(n286), .Z(n1803) );
  OAI21_X4 U1154 ( .B1(n2831), .B2(n360), .A(n2253), .ZN(n2219) );
  AOI222_X2 U1155 ( .A1(n3141), .A2(n421), .B1(n329), .B2(n418), .C1(n384), 
        .C2(n415), .ZN(n2253) );
  XOR2_X2 U1156 ( .A(n2220), .B(n286), .Z(n1804) );
  OAI21_X4 U1157 ( .B1(n2832), .B2(n360), .A(n2254), .ZN(n2220) );
  AOI222_X2 U1158 ( .A1(n3141), .A2(n418), .B1(n329), .B2(n415), .C1(n384), 
        .C2(n412), .ZN(n2254) );
  XOR2_X2 U1159 ( .A(n2221), .B(n286), .Z(n1805) );
  OAI21_X4 U1160 ( .B1(n2833), .B2(n360), .A(n2255), .ZN(n2221) );
  AOI222_X2 U1161 ( .A1(n3141), .A2(n415), .B1(n329), .B2(n412), .C1(n384), 
        .C2(n409), .ZN(n2255) );
  XOR2_X2 U1162 ( .A(n2222), .B(n286), .Z(n1806) );
  AOI222_X2 U1164 ( .A1(n3141), .A2(n412), .B1(n329), .B2(n409), .C1(n384), 
        .C2(n406), .ZN(n2256) );
  XOR2_X2 U1165 ( .A(n2223), .B(n286), .Z(n1807) );
  OAI21_X4 U1166 ( .B1(n2835), .B2(n360), .A(n2257), .ZN(n2223) );
  AOI222_X2 U1167 ( .A1(n3141), .A2(n409), .B1(n329), .B2(n406), .C1(n384), 
        .C2(n403), .ZN(n2257) );
  XOR2_X2 U1168 ( .A(n2224), .B(n286), .Z(n1808) );
  OAI21_X4 U1169 ( .B1(n2836), .B2(n360), .A(n2258), .ZN(n2224) );
  AOI222_X2 U1170 ( .A1(n3141), .A2(n406), .B1(n329), .B2(n403), .C1(n384), 
        .C2(n400), .ZN(n2258) );
  XOR2_X2 U1171 ( .A(n2225), .B(n286), .Z(n1809) );
  OAI21_X4 U1172 ( .B1(n2837), .B2(n360), .A(n2259), .ZN(n2225) );
  AOI222_X2 U1173 ( .A1(n307), .A2(n403), .B1(n329), .B2(n400), .C1(n384), 
        .C2(n397), .ZN(n2259) );
  XOR2_X2 U1174 ( .A(n2226), .B(n286), .Z(n1810) );
  OAI21_X4 U1175 ( .B1(n2838), .B2(n360), .A(n2260), .ZN(n2226) );
  AOI222_X2 U1176 ( .A1(n307), .A2(n400), .B1(n329), .B2(n397), .C1(n384), 
        .C2(n393), .ZN(n2260) );
  XOR2_X2 U1177 ( .A(n2227), .B(n286), .Z(n1811) );
  OAI21_X4 U1178 ( .B1(n2839), .B2(n360), .A(n2261), .ZN(n2227) );
  AOI222_X2 U1179 ( .A1(n307), .A2(n397), .B1(n329), .B2(n393), .C1(n384), 
        .C2(n390), .ZN(n2261) );
  XOR2_X2 U1180 ( .A(n2228), .B(n286), .Z(n1812) );
  OAI21_X4 U1181 ( .B1(n2840), .B2(n360), .A(n2262), .ZN(n2228) );
  XOR2_X2 U1183 ( .A(n2229), .B(n286), .Z(n1813) );
  OAI21_X4 U1184 ( .B1(n2841), .B2(n360), .A(n2263), .ZN(n2229) );
  AND2_X4 U1186 ( .A1(n307), .A2(n390), .ZN(n1382) );
  XOR2_X2 U1188 ( .A(n2264), .B(n283), .Z(n1815) );
  OAI21_X4 U1189 ( .B1(n2808), .B2(n357), .A(n2298), .ZN(n2264) );
  NAND2_X4 U1190 ( .A1(n382), .A2(n484), .ZN(n2298) );
  XOR2_X2 U1191 ( .A(n2265), .B(n283), .Z(n1816) );
  OAI21_X4 U1192 ( .B1(n2809), .B2(n357), .A(n2299), .ZN(n2265) );
  AOI21_X4 U1193 ( .B1(n382), .B2(n481), .A(n1383), .ZN(n2299) );
  AND2_X4 U1194 ( .A1(n327), .A2(n484), .ZN(n1383) );
  XOR2_X2 U1195 ( .A(n2266), .B(n283), .Z(n1817) );
  OAI21_X4 U1196 ( .B1(n2810), .B2(n357), .A(n2300), .ZN(n2266) );
  AOI222_X2 U1197 ( .A1(n3140), .A2(n484), .B1(n327), .B2(n481), .C1(n382), 
        .C2(n478), .ZN(n2300) );
  XOR2_X2 U1198 ( .A(n2267), .B(n283), .Z(n1818) );
  OAI21_X4 U1199 ( .B1(n2811), .B2(n357), .A(n2301), .ZN(n2267) );
  AOI222_X2 U1200 ( .A1(n3139), .A2(n481), .B1(n327), .B2(n478), .C1(n382), 
        .C2(n475), .ZN(n2301) );
  XOR2_X2 U1201 ( .A(n2268), .B(n283), .Z(n1819) );
  OAI21_X4 U1202 ( .B1(n2812), .B2(n357), .A(n2302), .ZN(n2268) );
  AOI222_X2 U1203 ( .A1(n3140), .A2(n478), .B1(n327), .B2(n475), .C1(n382), 
        .C2(n472), .ZN(n2302) );
  XOR2_X2 U1204 ( .A(n2269), .B(n283), .Z(n1820) );
  OAI21_X4 U1205 ( .B1(n2813), .B2(n357), .A(n2303), .ZN(n2269) );
  AOI222_X2 U1206 ( .A1(n3139), .A2(n475), .B1(n327), .B2(n472), .C1(n382), 
        .C2(n469), .ZN(n2303) );
  XOR2_X2 U1207 ( .A(n2270), .B(n283), .Z(n1821) );
  OAI21_X4 U1208 ( .B1(n2814), .B2(n357), .A(n2304), .ZN(n2270) );
  AOI222_X2 U1209 ( .A1(n3140), .A2(n472), .B1(n327), .B2(n469), .C1(n382), 
        .C2(n466), .ZN(n2304) );
  XOR2_X2 U1210 ( .A(n2271), .B(n283), .Z(n1822) );
  OAI21_X4 U1211 ( .B1(n2815), .B2(n357), .A(n2305), .ZN(n2271) );
  AOI222_X2 U1212 ( .A1(n3139), .A2(n469), .B1(n327), .B2(n466), .C1(n382), 
        .C2(n463), .ZN(n2305) );
  XOR2_X2 U1213 ( .A(n2272), .B(n283), .Z(n1823) );
  OAI21_X4 U1214 ( .B1(n2816), .B2(n357), .A(n2306), .ZN(n2272) );
  AOI222_X2 U1215 ( .A1(n3140), .A2(n466), .B1(n327), .B2(n463), .C1(n382), 
        .C2(n460), .ZN(n2306) );
  XOR2_X2 U1216 ( .A(n2273), .B(n283), .Z(n1824) );
  OAI21_X4 U1217 ( .B1(n2817), .B2(n357), .A(n2307), .ZN(n2273) );
  AOI222_X2 U1218 ( .A1(n3139), .A2(n463), .B1(n327), .B2(n460), .C1(n382), 
        .C2(n457), .ZN(n2307) );
  XOR2_X2 U1219 ( .A(n2274), .B(n283), .Z(n1825) );
  OAI21_X4 U1220 ( .B1(n2818), .B2(n357), .A(n2308), .ZN(n2274) );
  AOI222_X2 U1221 ( .A1(n3140), .A2(n460), .B1(n327), .B2(n457), .C1(n382), 
        .C2(n454), .ZN(n2308) );
  XOR2_X2 U1222 ( .A(n2275), .B(n283), .Z(n1826) );
  OAI21_X4 U1223 ( .B1(n2819), .B2(n357), .A(n2309), .ZN(n2275) );
  AOI222_X2 U1224 ( .A1(n3139), .A2(n457), .B1(n327), .B2(n454), .C1(n382), 
        .C2(n451), .ZN(n2309) );
  XOR2_X2 U1225 ( .A(n2276), .B(n283), .Z(n1827) );
  OAI21_X4 U1226 ( .B1(n2820), .B2(n357), .A(n2310), .ZN(n2276) );
  AOI222_X2 U1227 ( .A1(n3140), .A2(n454), .B1(n327), .B2(n451), .C1(n382), 
        .C2(n448), .ZN(n2310) );
  XOR2_X2 U1228 ( .A(n2277), .B(n283), .Z(n1828) );
  OAI21_X4 U1229 ( .B1(n2821), .B2(n357), .A(n2311), .ZN(n2277) );
  AOI222_X2 U1230 ( .A1(n3139), .A2(n451), .B1(n327), .B2(n448), .C1(n382), 
        .C2(n445), .ZN(n2311) );
  XOR2_X2 U1231 ( .A(n2278), .B(n283), .Z(n1829) );
  OAI21_X4 U1232 ( .B1(n2822), .B2(n357), .A(n2312), .ZN(n2278) );
  AOI222_X2 U1233 ( .A1(n3140), .A2(n448), .B1(n327), .B2(n445), .C1(n382), 
        .C2(n442), .ZN(n2312) );
  XOR2_X2 U1234 ( .A(n2279), .B(n283), .Z(n1830) );
  OAI21_X4 U1235 ( .B1(n2823), .B2(n357), .A(n2313), .ZN(n2279) );
  AOI222_X2 U1236 ( .A1(n3139), .A2(n445), .B1(n327), .B2(n442), .C1(n382), 
        .C2(n439), .ZN(n2313) );
  XOR2_X2 U1237 ( .A(n2280), .B(n283), .Z(n1831) );
  OAI21_X4 U1238 ( .B1(n2824), .B2(n357), .A(n2314), .ZN(n2280) );
  AOI222_X2 U1239 ( .A1(n3140), .A2(n442), .B1(n327), .B2(n439), .C1(n382), 
        .C2(n436), .ZN(n2314) );
  XOR2_X2 U1240 ( .A(n2281), .B(n283), .Z(n1832) );
  OAI21_X4 U1241 ( .B1(n2825), .B2(n357), .A(n2315), .ZN(n2281) );
  AOI222_X2 U1242 ( .A1(n3139), .A2(n439), .B1(n327), .B2(n436), .C1(n382), 
        .C2(n433), .ZN(n2315) );
  XOR2_X2 U1243 ( .A(n2282), .B(n283), .Z(n1833) );
  OAI21_X4 U1244 ( .B1(n2826), .B2(n357), .A(n2316), .ZN(n2282) );
  AOI222_X2 U1245 ( .A1(n3140), .A2(n436), .B1(n327), .B2(n433), .C1(n382), 
        .C2(n430), .ZN(n2316) );
  XOR2_X2 U1246 ( .A(n2283), .B(n283), .Z(n1834) );
  OAI21_X4 U1247 ( .B1(n2827), .B2(n357), .A(n2317), .ZN(n2283) );
  AOI222_X2 U1248 ( .A1(n3139), .A2(n433), .B1(n327), .B2(n430), .C1(n382), 
        .C2(n427), .ZN(n2317) );
  XOR2_X2 U1249 ( .A(n2284), .B(n283), .Z(n1835) );
  OAI21_X4 U1250 ( .B1(n2828), .B2(n357), .A(n2318), .ZN(n2284) );
  AOI222_X2 U1251 ( .A1(n3140), .A2(n430), .B1(n327), .B2(n427), .C1(n382), 
        .C2(n424), .ZN(n2318) );
  XOR2_X2 U1252 ( .A(n2285), .B(n283), .Z(n1836) );
  OAI21_X4 U1253 ( .B1(n2829), .B2(n357), .A(n2319), .ZN(n2285) );
  AOI222_X2 U1254 ( .A1(n3140), .A2(n427), .B1(n327), .B2(n424), .C1(n382), 
        .C2(n421), .ZN(n2319) );
  XOR2_X2 U1255 ( .A(n2286), .B(n283), .Z(n1837) );
  OAI21_X4 U1256 ( .B1(n2830), .B2(n357), .A(n2320), .ZN(n2286) );
  AOI222_X2 U1257 ( .A1(n3139), .A2(n424), .B1(n327), .B2(n421), .C1(n382), 
        .C2(n418), .ZN(n2320) );
  XOR2_X2 U1258 ( .A(n2287), .B(n283), .Z(n1838) );
  OAI21_X4 U1259 ( .B1(n2831), .B2(n357), .A(n2321), .ZN(n2287) );
  AOI222_X2 U1260 ( .A1(n3139), .A2(n421), .B1(n327), .B2(n418), .C1(n382), 
        .C2(n415), .ZN(n2321) );
  XOR2_X2 U1261 ( .A(n2288), .B(n283), .Z(n1839) );
  OAI21_X4 U1262 ( .B1(n2832), .B2(n357), .A(n2322), .ZN(n2288) );
  AOI222_X2 U1263 ( .A1(n3139), .A2(n418), .B1(n327), .B2(n415), .C1(n382), 
        .C2(n412), .ZN(n2322) );
  XOR2_X2 U1264 ( .A(n2289), .B(n283), .Z(n1840) );
  OAI21_X4 U1265 ( .B1(n2833), .B2(n357), .A(n2323), .ZN(n2289) );
  AOI222_X2 U1266 ( .A1(n3140), .A2(n415), .B1(n327), .B2(n412), .C1(n382), 
        .C2(n409), .ZN(n2323) );
  XOR2_X2 U1267 ( .A(n2290), .B(n283), .Z(n1841) );
  AOI222_X2 U1269 ( .A1(n3140), .A2(n412), .B1(n327), .B2(n409), .C1(n382), 
        .C2(n406), .ZN(n2324) );
  XOR2_X2 U1270 ( .A(n2291), .B(n283), .Z(n1842) );
  OAI21_X4 U1271 ( .B1(n2835), .B2(n357), .A(n2325), .ZN(n2291) );
  AOI222_X2 U1272 ( .A1(n3140), .A2(n409), .B1(n327), .B2(n406), .C1(n382), 
        .C2(n403), .ZN(n2325) );
  XOR2_X2 U1273 ( .A(n2292), .B(n283), .Z(n1843) );
  OAI21_X4 U1274 ( .B1(n2836), .B2(n357), .A(n2326), .ZN(n2292) );
  AOI222_X2 U1275 ( .A1(n3139), .A2(n406), .B1(n327), .B2(n403), .C1(n382), 
        .C2(n400), .ZN(n2326) );
  XOR2_X2 U1276 ( .A(n2293), .B(n283), .Z(n1844) );
  OAI21_X4 U1277 ( .B1(n2837), .B2(n357), .A(n2327), .ZN(n2293) );
  AOI222_X2 U1278 ( .A1(n3139), .A2(n403), .B1(n327), .B2(n400), .C1(n382), 
        .C2(n397), .ZN(n2327) );
  XOR2_X2 U1279 ( .A(n2294), .B(n283), .Z(n1845) );
  OAI21_X4 U1280 ( .B1(n2838), .B2(n357), .A(n2328), .ZN(n2294) );
  AOI222_X2 U1281 ( .A1(n3140), .A2(n400), .B1(n327), .B2(n397), .C1(n382), 
        .C2(n393), .ZN(n2328) );
  XOR2_X2 U1282 ( .A(n2295), .B(n283), .Z(n1846) );
  OAI21_X4 U1283 ( .B1(n2839), .B2(n357), .A(n2329), .ZN(n2295) );
  AOI222_X2 U1284 ( .A1(n3139), .A2(n397), .B1(n327), .B2(n393), .C1(n382), 
        .C2(n390), .ZN(n2329) );
  XOR2_X2 U1285 ( .A(n2296), .B(n283), .Z(n1847) );
  OAI21_X4 U1286 ( .B1(n2840), .B2(n357), .A(n2330), .ZN(n2296) );
  XOR2_X2 U1288 ( .A(n2297), .B(n283), .Z(n1848) );
  OAI21_X4 U1289 ( .B1(n2841), .B2(n357), .A(n2331), .ZN(n2297) );
  AND2_X4 U1291 ( .A1(n3139), .A2(n390), .ZN(n1385) );
  XOR2_X2 U1293 ( .A(n2332), .B(n280), .Z(n1850) );
  OAI21_X4 U1294 ( .B1(n2808), .B2(n354), .A(n2366), .ZN(n2332) );
  NAND2_X4 U1295 ( .A1(n380), .A2(n484), .ZN(n2366) );
  XOR2_X2 U1296 ( .A(n2333), .B(n280), .Z(n1851) );
  OAI21_X4 U1297 ( .B1(n2809), .B2(n354), .A(n2367), .ZN(n2333) );
  AOI21_X4 U1298 ( .B1(n380), .B2(n481), .A(n1386), .ZN(n2367) );
  AND2_X4 U1299 ( .A1(n325), .A2(n484), .ZN(n1386) );
  XOR2_X2 U1300 ( .A(n2334), .B(n280), .Z(n1852) );
  OAI21_X4 U1301 ( .B1(n2810), .B2(n354), .A(n2368), .ZN(n2334) );
  AOI222_X2 U1302 ( .A1(n3137), .A2(n484), .B1(n325), .B2(n481), .C1(n380), 
        .C2(n478), .ZN(n2368) );
  XOR2_X2 U1303 ( .A(n2335), .B(n280), .Z(n1853) );
  OAI21_X4 U1304 ( .B1(n2811), .B2(n354), .A(n2369), .ZN(n2335) );
  AOI222_X2 U1305 ( .A1(n3136), .A2(n481), .B1(n325), .B2(n478), .C1(n380), 
        .C2(n475), .ZN(n2369) );
  XOR2_X2 U1306 ( .A(n2336), .B(n280), .Z(n1854) );
  OAI21_X4 U1307 ( .B1(n2812), .B2(n354), .A(n2370), .ZN(n2336) );
  AOI222_X2 U1308 ( .A1(n3137), .A2(n478), .B1(n325), .B2(n475), .C1(n380), 
        .C2(n472), .ZN(n2370) );
  XOR2_X2 U1309 ( .A(n2337), .B(n280), .Z(n1855) );
  OAI21_X4 U1310 ( .B1(n2813), .B2(n354), .A(n2371), .ZN(n2337) );
  AOI222_X2 U1311 ( .A1(n3136), .A2(n475), .B1(n325), .B2(n472), .C1(n380), 
        .C2(n469), .ZN(n2371) );
  XOR2_X2 U1312 ( .A(n2338), .B(n280), .Z(n1856) );
  OAI21_X4 U1313 ( .B1(n2814), .B2(n354), .A(n2372), .ZN(n2338) );
  AOI222_X2 U1314 ( .A1(n3137), .A2(n472), .B1(n325), .B2(n469), .C1(n380), 
        .C2(n466), .ZN(n2372) );
  XOR2_X2 U1315 ( .A(n2339), .B(n280), .Z(n1857) );
  OAI21_X4 U1316 ( .B1(n2815), .B2(n354), .A(n2373), .ZN(n2339) );
  AOI222_X2 U1317 ( .A1(n3136), .A2(n469), .B1(n325), .B2(n466), .C1(n380), 
        .C2(n463), .ZN(n2373) );
  XOR2_X2 U1318 ( .A(n2340), .B(n280), .Z(n1858) );
  OAI21_X4 U1319 ( .B1(n2816), .B2(n354), .A(n2374), .ZN(n2340) );
  AOI222_X2 U1320 ( .A1(n3137), .A2(n466), .B1(n325), .B2(n463), .C1(n380), 
        .C2(n460), .ZN(n2374) );
  XOR2_X2 U1321 ( .A(n2341), .B(n280), .Z(n1859) );
  OAI21_X4 U1322 ( .B1(n2817), .B2(n354), .A(n2375), .ZN(n2341) );
  AOI222_X2 U1323 ( .A1(n3136), .A2(n463), .B1(n325), .B2(n460), .C1(n380), 
        .C2(n457), .ZN(n2375) );
  XOR2_X2 U1324 ( .A(n2342), .B(n280), .Z(n1860) );
  OAI21_X4 U1325 ( .B1(n2818), .B2(n354), .A(n2376), .ZN(n2342) );
  AOI222_X2 U1326 ( .A1(n3137), .A2(n460), .B1(n325), .B2(n457), .C1(n380), 
        .C2(n454), .ZN(n2376) );
  XOR2_X2 U1327 ( .A(n2343), .B(n280), .Z(n1861) );
  OAI21_X4 U1328 ( .B1(n2819), .B2(n354), .A(n2377), .ZN(n2343) );
  AOI222_X2 U1329 ( .A1(n3136), .A2(n457), .B1(n325), .B2(n454), .C1(n380), 
        .C2(n451), .ZN(n2377) );
  XOR2_X2 U1330 ( .A(n2344), .B(n280), .Z(n1862) );
  OAI21_X4 U1331 ( .B1(n2820), .B2(n354), .A(n2378), .ZN(n2344) );
  AOI222_X2 U1332 ( .A1(n3137), .A2(n454), .B1(n325), .B2(n451), .C1(n380), 
        .C2(n448), .ZN(n2378) );
  XOR2_X2 U1333 ( .A(n2345), .B(n280), .Z(n1863) );
  OAI21_X4 U1334 ( .B1(n2821), .B2(n354), .A(n2379), .ZN(n2345) );
  AOI222_X2 U1335 ( .A1(n3136), .A2(n451), .B1(n325), .B2(n448), .C1(n380), 
        .C2(n445), .ZN(n2379) );
  XOR2_X2 U1336 ( .A(n2346), .B(n280), .Z(n1864) );
  OAI21_X4 U1337 ( .B1(n2822), .B2(n354), .A(n2380), .ZN(n2346) );
  AOI222_X2 U1338 ( .A1(n3137), .A2(n448), .B1(n325), .B2(n445), .C1(n380), 
        .C2(n442), .ZN(n2380) );
  XOR2_X2 U1339 ( .A(n2347), .B(n280), .Z(n1865) );
  OAI21_X4 U1340 ( .B1(n2823), .B2(n354), .A(n2381), .ZN(n2347) );
  AOI222_X2 U1341 ( .A1(n3136), .A2(n445), .B1(n325), .B2(n442), .C1(n380), 
        .C2(n439), .ZN(n2381) );
  XOR2_X2 U1342 ( .A(n2348), .B(n280), .Z(n1866) );
  OAI21_X4 U1343 ( .B1(n2824), .B2(n354), .A(n2382), .ZN(n2348) );
  AOI222_X2 U1344 ( .A1(n3137), .A2(n442), .B1(n325), .B2(n439), .C1(n380), 
        .C2(n436), .ZN(n2382) );
  XOR2_X2 U1345 ( .A(n2349), .B(n280), .Z(n1867) );
  OAI21_X4 U1346 ( .B1(n2825), .B2(n354), .A(n2383), .ZN(n2349) );
  AOI222_X2 U1347 ( .A1(n3136), .A2(n439), .B1(n325), .B2(n436), .C1(n380), 
        .C2(n433), .ZN(n2383) );
  XOR2_X2 U1348 ( .A(n2350), .B(n280), .Z(n1868) );
  OAI21_X4 U1349 ( .B1(n2826), .B2(n354), .A(n2384), .ZN(n2350) );
  AOI222_X2 U1350 ( .A1(n3137), .A2(n436), .B1(n325), .B2(n433), .C1(n380), 
        .C2(n430), .ZN(n2384) );
  XOR2_X2 U1351 ( .A(n2351), .B(n280), .Z(n1869) );
  OAI21_X4 U1352 ( .B1(n2827), .B2(n354), .A(n2385), .ZN(n2351) );
  AOI222_X2 U1353 ( .A1(n3136), .A2(n433), .B1(n325), .B2(n430), .C1(n380), 
        .C2(n427), .ZN(n2385) );
  XOR2_X2 U1354 ( .A(n2352), .B(n280), .Z(n1870) );
  OAI21_X4 U1355 ( .B1(n2828), .B2(n354), .A(n2386), .ZN(n2352) );
  AOI222_X2 U1356 ( .A1(n3136), .A2(n430), .B1(n325), .B2(n427), .C1(n380), 
        .C2(n424), .ZN(n2386) );
  XOR2_X2 U1357 ( .A(n2353), .B(n280), .Z(n1871) );
  OAI21_X4 U1358 ( .B1(n2829), .B2(n354), .A(n2387), .ZN(n2353) );
  AOI222_X2 U1359 ( .A1(n3137), .A2(n427), .B1(n325), .B2(n424), .C1(n380), 
        .C2(n421), .ZN(n2387) );
  XOR2_X2 U1360 ( .A(n2354), .B(n280), .Z(n1872) );
  OAI21_X4 U1361 ( .B1(n2830), .B2(n354), .A(n2388), .ZN(n2354) );
  AOI222_X2 U1362 ( .A1(n3137), .A2(n424), .B1(n325), .B2(n421), .C1(n380), 
        .C2(n418), .ZN(n2388) );
  XOR2_X2 U1363 ( .A(n2355), .B(n280), .Z(n1873) );
  OAI21_X4 U1364 ( .B1(n2831), .B2(n354), .A(n2389), .ZN(n2355) );
  AOI222_X2 U1365 ( .A1(n3136), .A2(n421), .B1(n325), .B2(n418), .C1(n380), 
        .C2(n415), .ZN(n2389) );
  XOR2_X2 U1366 ( .A(n2356), .B(n280), .Z(n1874) );
  OAI21_X4 U1367 ( .B1(n2832), .B2(n354), .A(n2390), .ZN(n2356) );
  AOI222_X2 U1368 ( .A1(n3136), .A2(n418), .B1(n325), .B2(n415), .C1(n380), 
        .C2(n412), .ZN(n2390) );
  XOR2_X2 U1369 ( .A(n2357), .B(n280), .Z(n1875) );
  OAI21_X4 U1370 ( .B1(n2833), .B2(n354), .A(n2391), .ZN(n2357) );
  AOI222_X2 U1371 ( .A1(n3137), .A2(n415), .B1(n325), .B2(n412), .C1(n380), 
        .C2(n409), .ZN(n2391) );
  XOR2_X2 U1372 ( .A(n2358), .B(n280), .Z(n1876) );
  AOI222_X2 U1374 ( .A1(n3137), .A2(n412), .B1(n325), .B2(n409), .C1(n380), 
        .C2(n406), .ZN(n2392) );
  XOR2_X2 U1375 ( .A(n2359), .B(n280), .Z(n1877) );
  OAI21_X4 U1376 ( .B1(n2835), .B2(n354), .A(n2393), .ZN(n2359) );
  AOI222_X2 U1377 ( .A1(n3137), .A2(n409), .B1(n325), .B2(n406), .C1(n380), 
        .C2(n403), .ZN(n2393) );
  XOR2_X2 U1378 ( .A(n2360), .B(n280), .Z(n1878) );
  OAI21_X4 U1379 ( .B1(n2836), .B2(n354), .A(n2394), .ZN(n2360) );
  AOI222_X2 U1380 ( .A1(n3136), .A2(n406), .B1(n325), .B2(n403), .C1(n380), 
        .C2(n400), .ZN(n2394) );
  XOR2_X2 U1381 ( .A(n2361), .B(n280), .Z(n1879) );
  OAI21_X4 U1382 ( .B1(n2837), .B2(n354), .A(n2395), .ZN(n2361) );
  AOI222_X2 U1383 ( .A1(n3136), .A2(n403), .B1(n325), .B2(n400), .C1(n380), 
        .C2(n397), .ZN(n2395) );
  XOR2_X2 U1384 ( .A(n2362), .B(n280), .Z(n1880) );
  OAI21_X4 U1385 ( .B1(n2838), .B2(n354), .A(n2396), .ZN(n2362) );
  AOI222_X2 U1386 ( .A1(n3137), .A2(n400), .B1(n325), .B2(n397), .C1(n380), 
        .C2(n393), .ZN(n2396) );
  XOR2_X2 U1387 ( .A(n2363), .B(n280), .Z(n1881) );
  OAI21_X4 U1388 ( .B1(n2839), .B2(n354), .A(n2397), .ZN(n2363) );
  AOI222_X2 U1389 ( .A1(n3136), .A2(n397), .B1(n325), .B2(n393), .C1(n380), 
        .C2(n390), .ZN(n2397) );
  XOR2_X2 U1390 ( .A(n2364), .B(n280), .Z(n1882) );
  OAI21_X4 U1391 ( .B1(n2840), .B2(n354), .A(n2398), .ZN(n2364) );
  XOR2_X2 U1393 ( .A(n2365), .B(n280), .Z(n1883) );
  OAI21_X4 U1394 ( .B1(n2841), .B2(n354), .A(n2399), .ZN(n2365) );
  AND2_X4 U1396 ( .A1(n3136), .A2(n390), .ZN(n1388) );
  XOR2_X2 U1398 ( .A(n2400), .B(n277), .Z(n1885) );
  OAI21_X4 U1399 ( .B1(n2808), .B2(n351), .A(n2434), .ZN(n2400) );
  NAND2_X4 U1400 ( .A1(n378), .A2(n484), .ZN(n2434) );
  XOR2_X2 U1401 ( .A(n2401), .B(n277), .Z(n1886) );
  OAI21_X4 U1402 ( .B1(n2809), .B2(n351), .A(n2435), .ZN(n2401) );
  AOI21_X4 U1403 ( .B1(n378), .B2(n481), .A(n1389), .ZN(n2435) );
  AND2_X4 U1404 ( .A1(n323), .A2(n484), .ZN(n1389) );
  XOR2_X2 U1405 ( .A(n2402), .B(n277), .Z(n1887) );
  OAI21_X4 U1406 ( .B1(n2810), .B2(n351), .A(n2436), .ZN(n2402) );
  AOI222_X2 U1407 ( .A1(n3134), .A2(n484), .B1(n323), .B2(n481), .C1(n378), 
        .C2(n478), .ZN(n2436) );
  XOR2_X2 U1408 ( .A(n2403), .B(n277), .Z(n1888) );
  OAI21_X4 U1409 ( .B1(n2811), .B2(n351), .A(n2437), .ZN(n2403) );
  AOI222_X2 U1410 ( .A1(n3133), .A2(n481), .B1(n323), .B2(n478), .C1(n378), 
        .C2(n475), .ZN(n2437) );
  XOR2_X2 U1411 ( .A(n2404), .B(n277), .Z(n1889) );
  OAI21_X4 U1412 ( .B1(n2812), .B2(n351), .A(n2438), .ZN(n2404) );
  AOI222_X2 U1413 ( .A1(n3134), .A2(n478), .B1(n323), .B2(n475), .C1(n378), 
        .C2(n472), .ZN(n2438) );
  XOR2_X2 U1414 ( .A(n2405), .B(n277), .Z(n1890) );
  OAI21_X4 U1415 ( .B1(n2813), .B2(n351), .A(n2439), .ZN(n2405) );
  AOI222_X2 U1416 ( .A1(n3133), .A2(n475), .B1(n323), .B2(n472), .C1(n378), 
        .C2(n469), .ZN(n2439) );
  XOR2_X2 U1417 ( .A(n2406), .B(n277), .Z(n1891) );
  OAI21_X4 U1418 ( .B1(n2814), .B2(n351), .A(n2440), .ZN(n2406) );
  AOI222_X2 U1419 ( .A1(n3134), .A2(n472), .B1(n323), .B2(n469), .C1(n378), 
        .C2(n466), .ZN(n2440) );
  XOR2_X2 U1420 ( .A(n2407), .B(n277), .Z(n1892) );
  OAI21_X4 U1421 ( .B1(n2815), .B2(n351), .A(n2441), .ZN(n2407) );
  AOI222_X2 U1422 ( .A1(n3133), .A2(n469), .B1(n323), .B2(n466), .C1(n378), 
        .C2(n463), .ZN(n2441) );
  XOR2_X2 U1423 ( .A(n2408), .B(n277), .Z(n1893) );
  OAI21_X4 U1424 ( .B1(n2816), .B2(n351), .A(n2442), .ZN(n2408) );
  AOI222_X2 U1425 ( .A1(n3134), .A2(n466), .B1(n323), .B2(n463), .C1(n378), 
        .C2(n460), .ZN(n2442) );
  XOR2_X2 U1426 ( .A(n2409), .B(n277), .Z(n1894) );
  OAI21_X4 U1427 ( .B1(n2817), .B2(n351), .A(n2443), .ZN(n2409) );
  AOI222_X2 U1428 ( .A1(n3133), .A2(n463), .B1(n323), .B2(n460), .C1(n378), 
        .C2(n457), .ZN(n2443) );
  XOR2_X2 U1429 ( .A(n2410), .B(n277), .Z(n1895) );
  OAI21_X4 U1430 ( .B1(n2818), .B2(n351), .A(n2444), .ZN(n2410) );
  AOI222_X2 U1431 ( .A1(n3134), .A2(n460), .B1(n323), .B2(n457), .C1(n378), 
        .C2(n454), .ZN(n2444) );
  XOR2_X2 U1432 ( .A(n2411), .B(n277), .Z(n1896) );
  OAI21_X4 U1433 ( .B1(n2819), .B2(n351), .A(n2445), .ZN(n2411) );
  AOI222_X2 U1434 ( .A1(n3133), .A2(n457), .B1(n323), .B2(n454), .C1(n378), 
        .C2(n451), .ZN(n2445) );
  XOR2_X2 U1435 ( .A(n2412), .B(n277), .Z(n1897) );
  OAI21_X4 U1436 ( .B1(n2820), .B2(n351), .A(n2446), .ZN(n2412) );
  AOI222_X2 U1437 ( .A1(n3133), .A2(n454), .B1(n323), .B2(n451), .C1(n378), 
        .C2(n448), .ZN(n2446) );
  XOR2_X2 U1438 ( .A(n2413), .B(n277), .Z(n1898) );
  OAI21_X4 U1439 ( .B1(n2821), .B2(n351), .A(n2447), .ZN(n2413) );
  AOI222_X2 U1440 ( .A1(n3134), .A2(n451), .B1(n323), .B2(n448), .C1(n378), 
        .C2(n445), .ZN(n2447) );
  XOR2_X2 U1441 ( .A(n2414), .B(n277), .Z(n1899) );
  OAI21_X4 U1442 ( .B1(n2822), .B2(n351), .A(n2448), .ZN(n2414) );
  AOI222_X2 U1443 ( .A1(n3134), .A2(n448), .B1(n323), .B2(n445), .C1(n378), 
        .C2(n442), .ZN(n2448) );
  XOR2_X2 U1444 ( .A(n2415), .B(n277), .Z(n1900) );
  OAI21_X4 U1445 ( .B1(n2823), .B2(n351), .A(n2449), .ZN(n2415) );
  AOI222_X2 U1446 ( .A1(n3134), .A2(n445), .B1(n323), .B2(n442), .C1(n378), 
        .C2(n439), .ZN(n2449) );
  XOR2_X2 U1447 ( .A(n2416), .B(n277), .Z(n1901) );
  OAI21_X4 U1448 ( .B1(n2824), .B2(n351), .A(n2450), .ZN(n2416) );
  AOI222_X2 U1449 ( .A1(n3133), .A2(n442), .B1(n323), .B2(n439), .C1(n378), 
        .C2(n436), .ZN(n2450) );
  XOR2_X2 U1450 ( .A(n2417), .B(n277), .Z(n1902) );
  OAI21_X4 U1451 ( .B1(n2825), .B2(n351), .A(n2451), .ZN(n2417) );
  AOI222_X2 U1452 ( .A1(n3133), .A2(n439), .B1(n323), .B2(n436), .C1(n378), 
        .C2(n433), .ZN(n2451) );
  XOR2_X2 U1453 ( .A(n2418), .B(n277), .Z(n1903) );
  OAI21_X4 U1454 ( .B1(n2826), .B2(n351), .A(n2452), .ZN(n2418) );
  AOI222_X2 U1455 ( .A1(n3133), .A2(n436), .B1(n323), .B2(n433), .C1(n378), 
        .C2(n430), .ZN(n2452) );
  XOR2_X2 U1456 ( .A(n2419), .B(n277), .Z(n1904) );
  OAI21_X4 U1457 ( .B1(n2827), .B2(n351), .A(n2453), .ZN(n2419) );
  AOI222_X2 U1458 ( .A1(n3134), .A2(n433), .B1(n323), .B2(n430), .C1(n378), 
        .C2(n427), .ZN(n2453) );
  XOR2_X2 U1459 ( .A(n2420), .B(n277), .Z(n1905) );
  OAI21_X4 U1460 ( .B1(n2828), .B2(n351), .A(n2454), .ZN(n2420) );
  AOI222_X2 U1461 ( .A1(n3134), .A2(n430), .B1(n323), .B2(n427), .C1(n378), 
        .C2(n424), .ZN(n2454) );
  XOR2_X2 U1462 ( .A(n2421), .B(n277), .Z(n1906) );
  OAI21_X4 U1463 ( .B1(n2829), .B2(n351), .A(n2455), .ZN(n2421) );
  AOI222_X2 U1464 ( .A1(n3133), .A2(n427), .B1(n323), .B2(n424), .C1(n378), 
        .C2(n421), .ZN(n2455) );
  XOR2_X2 U1465 ( .A(n2422), .B(n277), .Z(n1907) );
  OAI21_X4 U1466 ( .B1(n2830), .B2(n351), .A(n2456), .ZN(n2422) );
  AOI222_X2 U1467 ( .A1(n3133), .A2(n424), .B1(n323), .B2(n421), .C1(n378), 
        .C2(n418), .ZN(n2456) );
  XOR2_X2 U1468 ( .A(n2423), .B(n277), .Z(n1908) );
  OAI21_X4 U1469 ( .B1(n2831), .B2(n351), .A(n2457), .ZN(n2423) );
  AOI222_X2 U1470 ( .A1(n3134), .A2(n421), .B1(n323), .B2(n418), .C1(n378), 
        .C2(n415), .ZN(n2457) );
  XOR2_X2 U1471 ( .A(n2424), .B(n277), .Z(n1909) );
  OAI21_X4 U1472 ( .B1(n2832), .B2(n351), .A(n2458), .ZN(n2424) );
  AOI222_X2 U1473 ( .A1(n3133), .A2(n418), .B1(n323), .B2(n415), .C1(n378), 
        .C2(n412), .ZN(n2458) );
  XOR2_X2 U1474 ( .A(n2425), .B(n277), .Z(n1910) );
  OAI21_X4 U1475 ( .B1(n2833), .B2(n351), .A(n2459), .ZN(n2425) );
  AOI222_X2 U1476 ( .A1(n3134), .A2(n415), .B1(n323), .B2(n412), .C1(n378), 
        .C2(n409), .ZN(n2459) );
  XOR2_X2 U1477 ( .A(n2426), .B(n277), .Z(n1911) );
  AOI222_X2 U1479 ( .A1(n3134), .A2(n412), .B1(n323), .B2(n409), .C1(n378), 
        .C2(n406), .ZN(n2460) );
  XOR2_X2 U1480 ( .A(n2427), .B(n277), .Z(n1912) );
  OAI21_X4 U1481 ( .B1(n2835), .B2(n351), .A(n2461), .ZN(n2427) );
  AOI222_X2 U1482 ( .A1(n3134), .A2(n409), .B1(n323), .B2(n406), .C1(n378), 
        .C2(n403), .ZN(n2461) );
  XOR2_X2 U1483 ( .A(n2428), .B(n277), .Z(n1913) );
  OAI21_X4 U1484 ( .B1(n2836), .B2(n351), .A(n2462), .ZN(n2428) );
  AOI222_X2 U1485 ( .A1(n3133), .A2(n406), .B1(n323), .B2(n403), .C1(n378), 
        .C2(n400), .ZN(n2462) );
  XOR2_X2 U1486 ( .A(n2429), .B(n277), .Z(n1914) );
  OAI21_X4 U1487 ( .B1(n2837), .B2(n351), .A(n2463), .ZN(n2429) );
  AOI222_X2 U1488 ( .A1(n3133), .A2(n403), .B1(n323), .B2(n400), .C1(n378), 
        .C2(n397), .ZN(n2463) );
  XOR2_X2 U1489 ( .A(n2430), .B(n277), .Z(n1915) );
  OAI21_X4 U1490 ( .B1(n2838), .B2(n351), .A(n2464), .ZN(n2430) );
  AOI222_X2 U1491 ( .A1(n3134), .A2(n400), .B1(n323), .B2(n397), .C1(n378), 
        .C2(n393), .ZN(n2464) );
  XOR2_X2 U1492 ( .A(n2431), .B(n277), .Z(n1916) );
  OAI21_X4 U1493 ( .B1(n2839), .B2(n351), .A(n2465), .ZN(n2431) );
  AOI222_X2 U1494 ( .A1(n3133), .A2(n397), .B1(n323), .B2(n393), .C1(n378), 
        .C2(n390), .ZN(n2465) );
  XOR2_X2 U1495 ( .A(n2432), .B(n277), .Z(n1917) );
  OAI21_X4 U1496 ( .B1(n2840), .B2(n351), .A(n2466), .ZN(n2432) );
  XOR2_X2 U1498 ( .A(n2433), .B(n277), .Z(n1918) );
  OAI21_X4 U1499 ( .B1(n2841), .B2(n351), .A(n2467), .ZN(n2433) );
  AND2_X4 U1501 ( .A1(n3133), .A2(n390), .ZN(n1391) );
  XOR2_X2 U1503 ( .A(n2468), .B(n274), .Z(n1920) );
  OAI21_X4 U1504 ( .B1(n2808), .B2(n348), .A(n2502), .ZN(n2468) );
  NAND2_X4 U1505 ( .A1(n376), .A2(n484), .ZN(n2502) );
  XOR2_X2 U1506 ( .A(n2469), .B(n274), .Z(n1921) );
  OAI21_X4 U1507 ( .B1(n2809), .B2(n348), .A(n2503), .ZN(n2469) );
  AOI21_X4 U1508 ( .B1(n376), .B2(n481), .A(n1392), .ZN(n2503) );
  AND2_X4 U1509 ( .A1(n321), .A2(n484), .ZN(n1392) );
  XOR2_X2 U1510 ( .A(n2470), .B(n274), .Z(n1922) );
  OAI21_X4 U1511 ( .B1(n2810), .B2(n348), .A(n2504), .ZN(n2470) );
  AOI222_X2 U1512 ( .A1(n3166), .A2(n484), .B1(n321), .B2(n481), .C1(n376), 
        .C2(n478), .ZN(n2504) );
  XOR2_X2 U1513 ( .A(n2471), .B(n274), .Z(n1923) );
  OAI21_X4 U1514 ( .B1(n2811), .B2(n348), .A(n2505), .ZN(n2471) );
  AOI222_X2 U1515 ( .A1(n3166), .A2(n481), .B1(n321), .B2(n478), .C1(n376), 
        .C2(n475), .ZN(n2505) );
  XOR2_X2 U1516 ( .A(n2472), .B(n274), .Z(n1924) );
  OAI21_X4 U1517 ( .B1(n2812), .B2(n348), .A(n2506), .ZN(n2472) );
  AOI222_X2 U1518 ( .A1(n3166), .A2(n478), .B1(n321), .B2(n475), .C1(n376), 
        .C2(n472), .ZN(n2506) );
  XOR2_X2 U1519 ( .A(n2473), .B(n274), .Z(n1925) );
  OAI21_X4 U1520 ( .B1(n2813), .B2(n348), .A(n2507), .ZN(n2473) );
  AOI222_X2 U1521 ( .A1(n3166), .A2(n475), .B1(n321), .B2(n472), .C1(n376), 
        .C2(n469), .ZN(n2507) );
  XOR2_X2 U1522 ( .A(n2474), .B(n274), .Z(n1926) );
  OAI21_X4 U1523 ( .B1(n2814), .B2(n348), .A(n2508), .ZN(n2474) );
  AOI222_X2 U1524 ( .A1(n3166), .A2(n472), .B1(n321), .B2(n469), .C1(n376), 
        .C2(n466), .ZN(n2508) );
  XOR2_X2 U1525 ( .A(n2475), .B(n274), .Z(n1927) );
  OAI21_X4 U1526 ( .B1(n2815), .B2(n348), .A(n2509), .ZN(n2475) );
  AOI222_X2 U1527 ( .A1(n3166), .A2(n469), .B1(n321), .B2(n466), .C1(n376), 
        .C2(n463), .ZN(n2509) );
  XOR2_X2 U1528 ( .A(n2476), .B(n274), .Z(n1928) );
  OAI21_X4 U1529 ( .B1(n2816), .B2(n348), .A(n2510), .ZN(n2476) );
  AOI222_X2 U1530 ( .A1(n3166), .A2(n466), .B1(n321), .B2(n463), .C1(n376), 
        .C2(n460), .ZN(n2510) );
  XOR2_X2 U1531 ( .A(n2477), .B(n274), .Z(n1929) );
  OAI21_X4 U1532 ( .B1(n2817), .B2(n348), .A(n2511), .ZN(n2477) );
  AOI222_X2 U1533 ( .A1(n3166), .A2(n463), .B1(n321), .B2(n460), .C1(n376), 
        .C2(n457), .ZN(n2511) );
  XOR2_X2 U1534 ( .A(n2478), .B(n274), .Z(n1930) );
  OAI21_X4 U1535 ( .B1(n2818), .B2(n348), .A(n2512), .ZN(n2478) );
  AOI222_X2 U1536 ( .A1(n3166), .A2(n460), .B1(n321), .B2(n457), .C1(n376), 
        .C2(n454), .ZN(n2512) );
  XOR2_X2 U1537 ( .A(n2479), .B(n274), .Z(n1931) );
  OAI21_X4 U1538 ( .B1(n2819), .B2(n348), .A(n2513), .ZN(n2479) );
  AOI222_X2 U1539 ( .A1(n3166), .A2(n457), .B1(n321), .B2(n454), .C1(n376), 
        .C2(n451), .ZN(n2513) );
  XOR2_X2 U1540 ( .A(n2480), .B(n274), .Z(n1932) );
  OAI21_X4 U1541 ( .B1(n2820), .B2(n348), .A(n2514), .ZN(n2480) );
  AOI222_X2 U1542 ( .A1(n3166), .A2(n454), .B1(n321), .B2(n451), .C1(n376), 
        .C2(n448), .ZN(n2514) );
  XOR2_X2 U1543 ( .A(n2481), .B(n274), .Z(n1933) );
  OAI21_X4 U1544 ( .B1(n2821), .B2(n348), .A(n2515), .ZN(n2481) );
  AOI222_X2 U1545 ( .A1(n3166), .A2(n451), .B1(n321), .B2(n448), .C1(n376), 
        .C2(n445), .ZN(n2515) );
  XOR2_X2 U1546 ( .A(n2482), .B(n274), .Z(n1934) );
  OAI21_X4 U1547 ( .B1(n2822), .B2(n348), .A(n2516), .ZN(n2482) );
  AOI222_X2 U1548 ( .A1(n3166), .A2(n448), .B1(n321), .B2(n445), .C1(n376), 
        .C2(n442), .ZN(n2516) );
  XOR2_X2 U1549 ( .A(n2483), .B(n274), .Z(n1935) );
  OAI21_X4 U1550 ( .B1(n2823), .B2(n348), .A(n2517), .ZN(n2483) );
  AOI222_X2 U1551 ( .A1(n3166), .A2(n445), .B1(n321), .B2(n442), .C1(n376), 
        .C2(n439), .ZN(n2517) );
  XOR2_X2 U1552 ( .A(n2484), .B(n274), .Z(n1936) );
  OAI21_X4 U1553 ( .B1(n2824), .B2(n348), .A(n2518), .ZN(n2484) );
  AOI222_X2 U1554 ( .A1(n3166), .A2(n442), .B1(n321), .B2(n439), .C1(n376), 
        .C2(n436), .ZN(n2518) );
  XOR2_X2 U1555 ( .A(n2485), .B(n274), .Z(n1937) );
  OAI21_X4 U1556 ( .B1(n2825), .B2(n348), .A(n2519), .ZN(n2485) );
  AOI222_X2 U1557 ( .A1(n3166), .A2(n439), .B1(n321), .B2(n436), .C1(n376), 
        .C2(n433), .ZN(n2519) );
  XOR2_X2 U1558 ( .A(n2486), .B(n274), .Z(n1938) );
  OAI21_X4 U1559 ( .B1(n2826), .B2(n348), .A(n2520), .ZN(n2486) );
  AOI222_X2 U1560 ( .A1(n3166), .A2(n436), .B1(n321), .B2(n433), .C1(n376), 
        .C2(n430), .ZN(n2520) );
  XOR2_X2 U1561 ( .A(n2487), .B(n274), .Z(n1939) );
  OAI21_X4 U1562 ( .B1(n2827), .B2(n348), .A(n2521), .ZN(n2487) );
  AOI222_X2 U1563 ( .A1(n3166), .A2(n433), .B1(n321), .B2(n430), .C1(n376), 
        .C2(n427), .ZN(n2521) );
  XOR2_X2 U1564 ( .A(n2488), .B(n274), .Z(n1940) );
  OAI21_X4 U1565 ( .B1(n2828), .B2(n348), .A(n2522), .ZN(n2488) );
  AOI222_X2 U1566 ( .A1(n3166), .A2(n430), .B1(n321), .B2(n427), .C1(n376), 
        .C2(n424), .ZN(n2522) );
  XOR2_X2 U1567 ( .A(n2489), .B(n274), .Z(n1941) );
  OAI21_X4 U1568 ( .B1(n2829), .B2(n348), .A(n2523), .ZN(n2489) );
  AOI222_X2 U1569 ( .A1(n3166), .A2(n427), .B1(n321), .B2(n424), .C1(n376), 
        .C2(n421), .ZN(n2523) );
  XOR2_X2 U1570 ( .A(n2490), .B(n274), .Z(n1942) );
  OAI21_X4 U1571 ( .B1(n2830), .B2(n348), .A(n2524), .ZN(n2490) );
  AOI222_X2 U1572 ( .A1(n3166), .A2(n424), .B1(n321), .B2(n421), .C1(n376), 
        .C2(n418), .ZN(n2524) );
  XOR2_X2 U1573 ( .A(n2491), .B(n274), .Z(n1943) );
  OAI21_X4 U1574 ( .B1(n2831), .B2(n348), .A(n2525), .ZN(n2491) );
  AOI222_X2 U1575 ( .A1(n3166), .A2(n421), .B1(n321), .B2(n418), .C1(n376), 
        .C2(n415), .ZN(n2525) );
  XOR2_X2 U1576 ( .A(n2492), .B(n274), .Z(n1944) );
  OAI21_X4 U1577 ( .B1(n2832), .B2(n348), .A(n2526), .ZN(n2492) );
  AOI222_X2 U1578 ( .A1(n3166), .A2(n418), .B1(n321), .B2(n415), .C1(n376), 
        .C2(n412), .ZN(n2526) );
  XOR2_X2 U1579 ( .A(n2493), .B(n274), .Z(n1945) );
  OAI21_X4 U1580 ( .B1(n2833), .B2(n348), .A(n2527), .ZN(n2493) );
  AOI222_X2 U1581 ( .A1(n3166), .A2(n415), .B1(n321), .B2(n412), .C1(n376), 
        .C2(n409), .ZN(n2527) );
  XOR2_X2 U1582 ( .A(n2494), .B(n274), .Z(n1946) );
  AOI222_X2 U1584 ( .A1(n3166), .A2(n412), .B1(n321), .B2(n409), .C1(n376), 
        .C2(n406), .ZN(n2528) );
  XOR2_X2 U1585 ( .A(n2495), .B(n274), .Z(n1947) );
  OAI21_X4 U1586 ( .B1(n2835), .B2(n348), .A(n2529), .ZN(n2495) );
  AOI222_X2 U1587 ( .A1(n3166), .A2(n409), .B1(n321), .B2(n406), .C1(n376), 
        .C2(n403), .ZN(n2529) );
  XOR2_X2 U1588 ( .A(n2496), .B(n274), .Z(n1948) );
  OAI21_X4 U1589 ( .B1(n2836), .B2(n348), .A(n2530), .ZN(n2496) );
  AOI222_X2 U1590 ( .A1(n3166), .A2(n406), .B1(n321), .B2(n403), .C1(n376), 
        .C2(n400), .ZN(n2530) );
  XOR2_X2 U1591 ( .A(n2497), .B(n274), .Z(n1949) );
  OAI21_X4 U1592 ( .B1(n2837), .B2(n348), .A(n2531), .ZN(n2497) );
  AOI222_X2 U1593 ( .A1(n3166), .A2(n403), .B1(n321), .B2(n400), .C1(n376), 
        .C2(n397), .ZN(n2531) );
  XOR2_X2 U1594 ( .A(n2498), .B(n274), .Z(n1950) );
  OAI21_X4 U1595 ( .B1(n2838), .B2(n348), .A(n2532), .ZN(n2498) );
  AOI222_X2 U1596 ( .A1(n3166), .A2(n400), .B1(n321), .B2(n397), .C1(n376), 
        .C2(n393), .ZN(n2532) );
  XOR2_X2 U1597 ( .A(n2499), .B(n274), .Z(n1951) );
  OAI21_X4 U1598 ( .B1(n2839), .B2(n348), .A(n2533), .ZN(n2499) );
  AOI222_X2 U1599 ( .A1(n3166), .A2(n397), .B1(n321), .B2(n393), .C1(n376), 
        .C2(n390), .ZN(n2533) );
  XOR2_X2 U1600 ( .A(n2500), .B(n274), .Z(n1952) );
  OAI21_X4 U1601 ( .B1(n2840), .B2(n348), .A(n2534), .ZN(n2500) );
  XOR2_X2 U1603 ( .A(n2501), .B(n274), .Z(n1953) );
  OAI21_X4 U1604 ( .B1(n2841), .B2(n348), .A(n2535), .ZN(n2501) );
  AND2_X4 U1606 ( .A1(n3166), .A2(n390), .ZN(n1394) );
  XOR2_X2 U1608 ( .A(n2536), .B(n271), .Z(n1955) );
  OAI21_X4 U1609 ( .B1(n2808), .B2(n345), .A(n2570), .ZN(n2536) );
  NAND2_X4 U1610 ( .A1(n374), .A2(n484), .ZN(n2570) );
  XOR2_X2 U1611 ( .A(n2537), .B(n271), .Z(n1956) );
  OAI21_X4 U1612 ( .B1(n2809), .B2(n345), .A(n2571), .ZN(n2537) );
  AOI21_X4 U1613 ( .B1(n374), .B2(n481), .A(n1395), .ZN(n2571) );
  AND2_X4 U1614 ( .A1(n319), .A2(n484), .ZN(n1395) );
  XOR2_X2 U1615 ( .A(n2538), .B(n271), .Z(n1957) );
  OAI21_X4 U1616 ( .B1(n2810), .B2(n345), .A(n2572), .ZN(n2538) );
  AOI222_X2 U1617 ( .A1(n297), .A2(n484), .B1(n319), .B2(n481), .C1(n374), 
        .C2(n478), .ZN(n2572) );
  XOR2_X2 U1618 ( .A(n2539), .B(n271), .Z(n1958) );
  OAI21_X4 U1619 ( .B1(n2811), .B2(n345), .A(n2573), .ZN(n2539) );
  AOI222_X2 U1620 ( .A1(n297), .A2(n481), .B1(n319), .B2(n478), .C1(n374), 
        .C2(n475), .ZN(n2573) );
  XOR2_X2 U1621 ( .A(n2540), .B(n271), .Z(n1959) );
  OAI21_X4 U1622 ( .B1(n2812), .B2(n345), .A(n2574), .ZN(n2540) );
  AOI222_X2 U1623 ( .A1(n297), .A2(n478), .B1(n319), .B2(n475), .C1(n374), 
        .C2(n472), .ZN(n2574) );
  XOR2_X2 U1624 ( .A(n2541), .B(n271), .Z(n1960) );
  OAI21_X4 U1625 ( .B1(n2813), .B2(n345), .A(n2575), .ZN(n2541) );
  AOI222_X2 U1626 ( .A1(n297), .A2(n475), .B1(n319), .B2(n472), .C1(n374), 
        .C2(n469), .ZN(n2575) );
  XOR2_X2 U1627 ( .A(n2542), .B(n271), .Z(n1961) );
  OAI21_X4 U1628 ( .B1(n2814), .B2(n345), .A(n2576), .ZN(n2542) );
  AOI222_X2 U1629 ( .A1(n297), .A2(n472), .B1(n319), .B2(n469), .C1(n374), 
        .C2(n466), .ZN(n2576) );
  XOR2_X2 U1630 ( .A(n2543), .B(n271), .Z(n1962) );
  OAI21_X4 U1631 ( .B1(n2815), .B2(n345), .A(n2577), .ZN(n2543) );
  AOI222_X2 U1632 ( .A1(n297), .A2(n469), .B1(n319), .B2(n466), .C1(n374), 
        .C2(n463), .ZN(n2577) );
  XOR2_X2 U1633 ( .A(n2544), .B(n271), .Z(n1963) );
  OAI21_X4 U1634 ( .B1(n2816), .B2(n345), .A(n2578), .ZN(n2544) );
  AOI222_X2 U1635 ( .A1(n297), .A2(n466), .B1(n319), .B2(n463), .C1(n374), 
        .C2(n460), .ZN(n2578) );
  XOR2_X2 U1636 ( .A(n2545), .B(n271), .Z(n1964) );
  OAI21_X4 U1637 ( .B1(n2817), .B2(n345), .A(n2579), .ZN(n2545) );
  AOI222_X2 U1638 ( .A1(n297), .A2(n463), .B1(n319), .B2(n460), .C1(n374), 
        .C2(n457), .ZN(n2579) );
  XOR2_X2 U1639 ( .A(n2546), .B(n271), .Z(n1965) );
  OAI21_X4 U1640 ( .B1(n2818), .B2(n345), .A(n2580), .ZN(n2546) );
  AOI222_X2 U1641 ( .A1(n297), .A2(n460), .B1(n319), .B2(n457), .C1(n374), 
        .C2(n454), .ZN(n2580) );
  XOR2_X2 U1642 ( .A(n2547), .B(n271), .Z(n1966) );
  OAI21_X4 U1643 ( .B1(n2819), .B2(n345), .A(n2581), .ZN(n2547) );
  AOI222_X2 U1644 ( .A1(n297), .A2(n457), .B1(n319), .B2(n454), .C1(n374), 
        .C2(n451), .ZN(n2581) );
  XOR2_X2 U1645 ( .A(n2548), .B(n271), .Z(n1967) );
  OAI21_X4 U1646 ( .B1(n2820), .B2(n345), .A(n2582), .ZN(n2548) );
  AOI222_X2 U1647 ( .A1(n297), .A2(n454), .B1(n319), .B2(n451), .C1(n374), 
        .C2(n448), .ZN(n2582) );
  XOR2_X2 U1648 ( .A(n2549), .B(n271), .Z(n1968) );
  OAI21_X4 U1649 ( .B1(n2821), .B2(n345), .A(n2583), .ZN(n2549) );
  AOI222_X2 U1650 ( .A1(n297), .A2(n451), .B1(n319), .B2(n448), .C1(n374), 
        .C2(n445), .ZN(n2583) );
  XOR2_X2 U1651 ( .A(n2550), .B(n271), .Z(n1969) );
  OAI21_X4 U1652 ( .B1(n2822), .B2(n345), .A(n2584), .ZN(n2550) );
  AOI222_X2 U1653 ( .A1(n297), .A2(n448), .B1(n319), .B2(n445), .C1(n374), 
        .C2(n442), .ZN(n2584) );
  XOR2_X2 U1654 ( .A(n2551), .B(n271), .Z(n1970) );
  OAI21_X4 U1655 ( .B1(n2823), .B2(n345), .A(n2585), .ZN(n2551) );
  AOI222_X2 U1656 ( .A1(n297), .A2(n445), .B1(n319), .B2(n442), .C1(n374), 
        .C2(n439), .ZN(n2585) );
  XOR2_X2 U1657 ( .A(n2552), .B(n271), .Z(n1971) );
  OAI21_X4 U1658 ( .B1(n2824), .B2(n345), .A(n2586), .ZN(n2552) );
  AOI222_X2 U1659 ( .A1(n297), .A2(n442), .B1(n319), .B2(n439), .C1(n374), 
        .C2(n436), .ZN(n2586) );
  XOR2_X2 U1660 ( .A(n2553), .B(n271), .Z(n1972) );
  OAI21_X4 U1661 ( .B1(n2825), .B2(n345), .A(n2587), .ZN(n2553) );
  AOI222_X2 U1662 ( .A1(n297), .A2(n439), .B1(n319), .B2(n436), .C1(n374), 
        .C2(n433), .ZN(n2587) );
  XOR2_X2 U1663 ( .A(n2554), .B(n271), .Z(n1973) );
  OAI21_X4 U1664 ( .B1(n2826), .B2(n345), .A(n2588), .ZN(n2554) );
  AOI222_X2 U1665 ( .A1(n297), .A2(n436), .B1(n319), .B2(n433), .C1(n374), 
        .C2(n430), .ZN(n2588) );
  XOR2_X2 U1666 ( .A(n2555), .B(n271), .Z(n1974) );
  OAI21_X4 U1667 ( .B1(n2827), .B2(n345), .A(n2589), .ZN(n2555) );
  AOI222_X2 U1668 ( .A1(n297), .A2(n433), .B1(n319), .B2(n430), .C1(n374), 
        .C2(n427), .ZN(n2589) );
  XOR2_X2 U1669 ( .A(n2556), .B(n271), .Z(n1975) );
  OAI21_X4 U1670 ( .B1(n2828), .B2(n345), .A(n2590), .ZN(n2556) );
  AOI222_X2 U1671 ( .A1(n297), .A2(n430), .B1(n319), .B2(n427), .C1(n374), 
        .C2(n424), .ZN(n2590) );
  XOR2_X2 U1672 ( .A(n2557), .B(n271), .Z(n1976) );
  OAI21_X4 U1673 ( .B1(n2829), .B2(n345), .A(n2591), .ZN(n2557) );
  AOI222_X2 U1674 ( .A1(n297), .A2(n427), .B1(n319), .B2(n424), .C1(n374), 
        .C2(n421), .ZN(n2591) );
  XOR2_X2 U1675 ( .A(n2558), .B(n271), .Z(n1977) );
  OAI21_X4 U1676 ( .B1(n2830), .B2(n345), .A(n2592), .ZN(n2558) );
  AOI222_X2 U1677 ( .A1(n297), .A2(n424), .B1(n319), .B2(n421), .C1(n374), 
        .C2(n418), .ZN(n2592) );
  XOR2_X2 U1678 ( .A(n2559), .B(n271), .Z(n1978) );
  OAI21_X4 U1679 ( .B1(n2831), .B2(n345), .A(n2593), .ZN(n2559) );
  AOI222_X2 U1680 ( .A1(n297), .A2(n421), .B1(n319), .B2(n418), .C1(n374), 
        .C2(n415), .ZN(n2593) );
  XOR2_X2 U1681 ( .A(n2560), .B(n271), .Z(n1979) );
  OAI21_X4 U1682 ( .B1(n2832), .B2(n345), .A(n2594), .ZN(n2560) );
  AOI222_X2 U1683 ( .A1(n297), .A2(n418), .B1(n319), .B2(n415), .C1(n374), 
        .C2(n412), .ZN(n2594) );
  XOR2_X2 U1684 ( .A(n2561), .B(n271), .Z(n1980) );
  OAI21_X4 U1685 ( .B1(n2833), .B2(n345), .A(n2595), .ZN(n2561) );
  AOI222_X2 U1686 ( .A1(n297), .A2(n415), .B1(n319), .B2(n412), .C1(n374), 
        .C2(n409), .ZN(n2595) );
  XOR2_X2 U1687 ( .A(n2562), .B(n271), .Z(n1981) );
  AOI222_X2 U1689 ( .A1(n297), .A2(n412), .B1(n319), .B2(n409), .C1(n374), 
        .C2(n406), .ZN(n2596) );
  XOR2_X2 U1690 ( .A(n2563), .B(n271), .Z(n1982) );
  OAI21_X4 U1691 ( .B1(n2835), .B2(n345), .A(n2597), .ZN(n2563) );
  AOI222_X2 U1692 ( .A1(n297), .A2(n409), .B1(n319), .B2(n406), .C1(n374), 
        .C2(n403), .ZN(n2597) );
  XOR2_X2 U1693 ( .A(n2564), .B(n271), .Z(n1983) );
  OAI21_X4 U1694 ( .B1(n2836), .B2(n345), .A(n2598), .ZN(n2564) );
  AOI222_X2 U1695 ( .A1(n297), .A2(n406), .B1(n319), .B2(n403), .C1(n374), 
        .C2(n400), .ZN(n2598) );
  XOR2_X2 U1696 ( .A(n2565), .B(n271), .Z(n1984) );
  OAI21_X4 U1697 ( .B1(n2837), .B2(n345), .A(n2599), .ZN(n2565) );
  AOI222_X2 U1698 ( .A1(n297), .A2(n403), .B1(n319), .B2(n400), .C1(n374), 
        .C2(n397), .ZN(n2599) );
  XOR2_X2 U1699 ( .A(n2566), .B(n271), .Z(n1985) );
  OAI21_X4 U1700 ( .B1(n2838), .B2(n345), .A(n2600), .ZN(n2566) );
  AOI222_X2 U1701 ( .A1(n297), .A2(n400), .B1(n319), .B2(n397), .C1(n374), 
        .C2(n393), .ZN(n2600) );
  XOR2_X2 U1702 ( .A(n2567), .B(n271), .Z(n1986) );
  OAI21_X4 U1703 ( .B1(n2839), .B2(n345), .A(n2601), .ZN(n2567) );
  AOI222_X2 U1704 ( .A1(n297), .A2(n397), .B1(n319), .B2(n393), .C1(n374), 
        .C2(n390), .ZN(n2601) );
  XOR2_X2 U1705 ( .A(n2568), .B(n271), .Z(n1987) );
  OAI21_X4 U1706 ( .B1(n2840), .B2(n345), .A(n2602), .ZN(n2568) );
  AND2_X4 U1711 ( .A1(n297), .A2(n390), .ZN(n1397) );
  XOR2_X2 U1713 ( .A(n2604), .B(n268), .Z(n1990) );
  OAI21_X4 U1714 ( .B1(n2808), .B2(n342), .A(n2638), .ZN(n2604) );
  NAND2_X4 U1715 ( .A1(n3169), .A2(n484), .ZN(n2638) );
  XOR2_X2 U1716 ( .A(n2605), .B(n268), .Z(n1991) );
  OAI21_X4 U1717 ( .B1(n2809), .B2(n342), .A(n2639), .ZN(n2605) );
  AOI21_X4 U1718 ( .B1(n3169), .B2(n481), .A(n1398), .ZN(n2639) );
  AND2_X4 U1719 ( .A1(n317), .A2(n484), .ZN(n1398) );
  XOR2_X2 U1720 ( .A(n2606), .B(n268), .Z(n1992) );
  OAI21_X4 U1721 ( .B1(n2810), .B2(n342), .A(n2640), .ZN(n2606) );
  AOI222_X2 U1722 ( .A1(n295), .A2(n484), .B1(n317), .B2(n481), .C1(n3169), 
        .C2(n478), .ZN(n2640) );
  XOR2_X2 U1723 ( .A(n2607), .B(n268), .Z(n1993) );
  OAI21_X4 U1724 ( .B1(n2811), .B2(n342), .A(n2641), .ZN(n2607) );
  AOI222_X2 U1725 ( .A1(n295), .A2(n481), .B1(n317), .B2(n478), .C1(n3169), 
        .C2(n475), .ZN(n2641) );
  XOR2_X2 U1726 ( .A(n2608), .B(n268), .Z(n1994) );
  OAI21_X4 U1727 ( .B1(n2812), .B2(n342), .A(n2642), .ZN(n2608) );
  AOI222_X2 U1728 ( .A1(n295), .A2(n478), .B1(n317), .B2(n475), .C1(n3169), 
        .C2(n472), .ZN(n2642) );
  XOR2_X2 U1729 ( .A(n2609), .B(n268), .Z(n1995) );
  OAI21_X4 U1730 ( .B1(n2813), .B2(n342), .A(n2643), .ZN(n2609) );
  AOI222_X2 U1731 ( .A1(n295), .A2(n475), .B1(n317), .B2(n472), .C1(n3169), 
        .C2(n469), .ZN(n2643) );
  XOR2_X2 U1732 ( .A(n2610), .B(n268), .Z(n1996) );
  OAI21_X4 U1733 ( .B1(n2814), .B2(n342), .A(n2644), .ZN(n2610) );
  AOI222_X2 U1734 ( .A1(n295), .A2(n472), .B1(n317), .B2(n469), .C1(n3169), 
        .C2(n466), .ZN(n2644) );
  XOR2_X2 U1735 ( .A(n2611), .B(n268), .Z(n1997) );
  OAI21_X4 U1736 ( .B1(n2815), .B2(n342), .A(n2645), .ZN(n2611) );
  AOI222_X2 U1737 ( .A1(n295), .A2(n469), .B1(n317), .B2(n466), .C1(n3169), 
        .C2(n463), .ZN(n2645) );
  XOR2_X2 U1738 ( .A(n2612), .B(n268), .Z(n1998) );
  OAI21_X4 U1739 ( .B1(n2816), .B2(n342), .A(n2646), .ZN(n2612) );
  AOI222_X2 U1740 ( .A1(n295), .A2(n466), .B1(n317), .B2(n463), .C1(n3169), 
        .C2(n460), .ZN(n2646) );
  XOR2_X2 U1741 ( .A(n2613), .B(n268), .Z(n1999) );
  OAI21_X4 U1742 ( .B1(n2817), .B2(n342), .A(n2647), .ZN(n2613) );
  AOI222_X2 U1743 ( .A1(n295), .A2(n463), .B1(n317), .B2(n460), .C1(n3169), 
        .C2(n457), .ZN(n2647) );
  XOR2_X2 U1744 ( .A(n2614), .B(n268), .Z(n2000) );
  OAI21_X4 U1745 ( .B1(n2818), .B2(n342), .A(n2648), .ZN(n2614) );
  AOI222_X2 U1746 ( .A1(n295), .A2(n460), .B1(n317), .B2(n457), .C1(n3169), 
        .C2(n454), .ZN(n2648) );
  XOR2_X2 U1747 ( .A(n2615), .B(n268), .Z(n2001) );
  OAI21_X4 U1748 ( .B1(n2819), .B2(n342), .A(n2649), .ZN(n2615) );
  AOI222_X2 U1749 ( .A1(n295), .A2(n457), .B1(n317), .B2(n454), .C1(n3169), 
        .C2(n451), .ZN(n2649) );
  XOR2_X2 U1750 ( .A(n2616), .B(n268), .Z(n2002) );
  OAI21_X4 U1751 ( .B1(n2820), .B2(n342), .A(n2650), .ZN(n2616) );
  AOI222_X2 U1752 ( .A1(n295), .A2(n454), .B1(n317), .B2(n451), .C1(n3169), 
        .C2(n448), .ZN(n2650) );
  XOR2_X2 U1753 ( .A(n2617), .B(n268), .Z(n2003) );
  OAI21_X4 U1754 ( .B1(n2821), .B2(n342), .A(n2651), .ZN(n2617) );
  AOI222_X2 U1755 ( .A1(n295), .A2(n451), .B1(n317), .B2(n448), .C1(n3169), 
        .C2(n445), .ZN(n2651) );
  XOR2_X2 U1756 ( .A(n2618), .B(n268), .Z(n2004) );
  OAI21_X4 U1757 ( .B1(n2822), .B2(n342), .A(n2652), .ZN(n2618) );
  AOI222_X2 U1758 ( .A1(n295), .A2(n448), .B1(n317), .B2(n445), .C1(n3169), 
        .C2(n442), .ZN(n2652) );
  XOR2_X2 U1759 ( .A(n2619), .B(n268), .Z(n2005) );
  OAI21_X4 U1760 ( .B1(n2823), .B2(n342), .A(n2653), .ZN(n2619) );
  AOI222_X2 U1761 ( .A1(n295), .A2(n445), .B1(n317), .B2(n442), .C1(n3169), 
        .C2(n439), .ZN(n2653) );
  XOR2_X2 U1762 ( .A(n2620), .B(n268), .Z(n2006) );
  OAI21_X4 U1763 ( .B1(n2824), .B2(n342), .A(n2654), .ZN(n2620) );
  AOI222_X2 U1764 ( .A1(n295), .A2(n442), .B1(n317), .B2(n439), .C1(n3169), 
        .C2(n436), .ZN(n2654) );
  XOR2_X2 U1765 ( .A(n2621), .B(n268), .Z(n2007) );
  OAI21_X4 U1766 ( .B1(n2825), .B2(n342), .A(n2655), .ZN(n2621) );
  AOI222_X2 U1767 ( .A1(n295), .A2(n439), .B1(n317), .B2(n436), .C1(n3169), 
        .C2(n433), .ZN(n2655) );
  XOR2_X2 U1768 ( .A(n2622), .B(n268), .Z(n2008) );
  OAI21_X4 U1769 ( .B1(n2826), .B2(n342), .A(n2656), .ZN(n2622) );
  AOI222_X2 U1770 ( .A1(n295), .A2(n436), .B1(n317), .B2(n433), .C1(n3169), 
        .C2(n430), .ZN(n2656) );
  XOR2_X2 U1771 ( .A(n2623), .B(n268), .Z(n2009) );
  OAI21_X4 U1772 ( .B1(n2827), .B2(n342), .A(n2657), .ZN(n2623) );
  AOI222_X2 U1773 ( .A1(n295), .A2(n433), .B1(n317), .B2(n430), .C1(n3169), 
        .C2(n427), .ZN(n2657) );
  XOR2_X2 U1774 ( .A(n2624), .B(n268), .Z(n2010) );
  OAI21_X4 U1775 ( .B1(n2828), .B2(n342), .A(n2658), .ZN(n2624) );
  AOI222_X2 U1776 ( .A1(n295), .A2(n430), .B1(n317), .B2(n427), .C1(n3169), 
        .C2(n424), .ZN(n2658) );
  XOR2_X2 U1777 ( .A(n2625), .B(n268), .Z(n2011) );
  OAI21_X4 U1778 ( .B1(n2829), .B2(n342), .A(n2659), .ZN(n2625) );
  AOI222_X2 U1779 ( .A1(n295), .A2(n427), .B1(n317), .B2(n424), .C1(n3169), 
        .C2(n421), .ZN(n2659) );
  XOR2_X2 U1780 ( .A(n2626), .B(n268), .Z(n2012) );
  OAI21_X4 U1781 ( .B1(n2830), .B2(n342), .A(n2660), .ZN(n2626) );
  AOI222_X2 U1782 ( .A1(n295), .A2(n424), .B1(n317), .B2(n421), .C1(n3169), 
        .C2(n418), .ZN(n2660) );
  XOR2_X2 U1783 ( .A(n2627), .B(n268), .Z(n2013) );
  OAI21_X4 U1784 ( .B1(n2831), .B2(n342), .A(n2661), .ZN(n2627) );
  AOI222_X2 U1785 ( .A1(n295), .A2(n421), .B1(n317), .B2(n418), .C1(n3169), 
        .C2(n415), .ZN(n2661) );
  XOR2_X2 U1786 ( .A(n2628), .B(n268), .Z(n2014) );
  OAI21_X4 U1787 ( .B1(n2832), .B2(n342), .A(n2662), .ZN(n2628) );
  AOI222_X2 U1788 ( .A1(n295), .A2(n418), .B1(n317), .B2(n415), .C1(n3169), 
        .C2(n412), .ZN(n2662) );
  XOR2_X2 U1789 ( .A(n2629), .B(n268), .Z(n2015) );
  OAI21_X4 U1790 ( .B1(n2833), .B2(n342), .A(n2663), .ZN(n2629) );
  AOI222_X2 U1791 ( .A1(n295), .A2(n415), .B1(n317), .B2(n412), .C1(n3169), 
        .C2(n409), .ZN(n2663) );
  XOR2_X2 U1792 ( .A(n2630), .B(n268), .Z(n2016) );
  AOI222_X2 U1794 ( .A1(n295), .A2(n412), .B1(n317), .B2(n409), .C1(n3169), 
        .C2(n406), .ZN(n2664) );
  XOR2_X2 U1795 ( .A(n2631), .B(n268), .Z(n2017) );
  OAI21_X4 U1796 ( .B1(n2835), .B2(n342), .A(n2665), .ZN(n2631) );
  AOI222_X2 U1797 ( .A1(n295), .A2(n409), .B1(n317), .B2(n406), .C1(n3169), 
        .C2(n403), .ZN(n2665) );
  XOR2_X2 U1798 ( .A(n2632), .B(n268), .Z(n2018) );
  OAI21_X4 U1799 ( .B1(n2836), .B2(n342), .A(n2666), .ZN(n2632) );
  AOI222_X2 U1800 ( .A1(n295), .A2(n406), .B1(n317), .B2(n403), .C1(n3169), 
        .C2(n400), .ZN(n2666) );
  XOR2_X2 U1801 ( .A(n2633), .B(n268), .Z(n2019) );
  OAI21_X4 U1802 ( .B1(n2837), .B2(n342), .A(n2667), .ZN(n2633) );
  AOI222_X2 U1803 ( .A1(n295), .A2(n403), .B1(n317), .B2(n400), .C1(n3169), 
        .C2(n397), .ZN(n2667) );
  XOR2_X2 U1804 ( .A(n2634), .B(n268), .Z(n2020) );
  OAI21_X4 U1805 ( .B1(n2838), .B2(n342), .A(n2668), .ZN(n2634) );
  AOI222_X2 U1806 ( .A1(n295), .A2(n400), .B1(n317), .B2(n397), .C1(n3169), 
        .C2(n393), .ZN(n2668) );
  XOR2_X2 U1807 ( .A(n2635), .B(n268), .Z(n2021) );
  OAI21_X4 U1808 ( .B1(n2839), .B2(n342), .A(n2669), .ZN(n2635) );
  AOI222_X2 U1809 ( .A1(n295), .A2(n397), .B1(n317), .B2(n393), .C1(n3168), 
        .C2(n390), .ZN(n2669) );
  XOR2_X2 U1810 ( .A(n2636), .B(n268), .Z(n2022) );
  AND2_X4 U1816 ( .A1(n295), .A2(n390), .ZN(n1400) );
  XOR2_X2 U1818 ( .A(n2672), .B(n265), .Z(n2025) );
  OAI21_X4 U1819 ( .B1(n2808), .B2(n339), .A(n2706), .ZN(n2672) );
  NAND2_X4 U1820 ( .A1(n370), .A2(n484), .ZN(n2706) );
  XOR2_X2 U1821 ( .A(n2673), .B(n265), .Z(n2026) );
  OAI21_X4 U1822 ( .B1(n2809), .B2(n339), .A(n2707), .ZN(n2673) );
  AOI21_X4 U1823 ( .B1(n370), .B2(n481), .A(n1401), .ZN(n2707) );
  AND2_X4 U1824 ( .A1(n315), .A2(n484), .ZN(n1401) );
  XOR2_X2 U1825 ( .A(n2674), .B(n265), .Z(n2027) );
  OAI21_X4 U1826 ( .B1(n2810), .B2(n339), .A(n2708), .ZN(n2674) );
  AOI222_X2 U1827 ( .A1(n3213), .A2(n484), .B1(n315), .B2(n481), .C1(n370), 
        .C2(n478), .ZN(n2708) );
  XOR2_X2 U1828 ( .A(n2675), .B(n265), .Z(n2028) );
  OAI21_X4 U1829 ( .B1(n2811), .B2(n339), .A(n2709), .ZN(n2675) );
  AOI222_X2 U1830 ( .A1(n3213), .A2(n481), .B1(n315), .B2(n478), .C1(n370), 
        .C2(n475), .ZN(n2709) );
  XOR2_X2 U1831 ( .A(n2676), .B(n265), .Z(n2029) );
  OAI21_X4 U1832 ( .B1(n2812), .B2(n339), .A(n2710), .ZN(n2676) );
  AOI222_X2 U1833 ( .A1(n3213), .A2(n478), .B1(n315), .B2(n475), .C1(n370), 
        .C2(n472), .ZN(n2710) );
  XOR2_X2 U1834 ( .A(n2677), .B(n265), .Z(n2030) );
  OAI21_X4 U1835 ( .B1(n2813), .B2(n339), .A(n2711), .ZN(n2677) );
  AOI222_X2 U1836 ( .A1(n3213), .A2(n475), .B1(n315), .B2(n472), .C1(n370), 
        .C2(n469), .ZN(n2711) );
  XOR2_X2 U1837 ( .A(n2678), .B(n265), .Z(n2031) );
  OAI21_X4 U1838 ( .B1(n2814), .B2(n339), .A(n2712), .ZN(n2678) );
  AOI222_X2 U1839 ( .A1(n3213), .A2(n472), .B1(n315), .B2(n469), .C1(n370), 
        .C2(n466), .ZN(n2712) );
  XOR2_X2 U1840 ( .A(n2679), .B(n265), .Z(n2032) );
  OAI21_X4 U1841 ( .B1(n2815), .B2(n339), .A(n2713), .ZN(n2679) );
  AOI222_X2 U1842 ( .A1(n3213), .A2(n469), .B1(n315), .B2(n466), .C1(n370), 
        .C2(n463), .ZN(n2713) );
  XOR2_X2 U1843 ( .A(n2680), .B(n265), .Z(n2033) );
  OAI21_X4 U1844 ( .B1(n2816), .B2(n339), .A(n2714), .ZN(n2680) );
  AOI222_X2 U1845 ( .A1(n3213), .A2(n466), .B1(n315), .B2(n463), .C1(n370), 
        .C2(n460), .ZN(n2714) );
  XOR2_X2 U1846 ( .A(n2681), .B(n265), .Z(n2034) );
  OAI21_X4 U1847 ( .B1(n2817), .B2(n339), .A(n2715), .ZN(n2681) );
  AOI222_X2 U1848 ( .A1(n3213), .A2(n463), .B1(n315), .B2(n460), .C1(n370), 
        .C2(n457), .ZN(n2715) );
  XOR2_X2 U1849 ( .A(n2682), .B(n265), .Z(n2035) );
  OAI21_X4 U1850 ( .B1(n2818), .B2(n339), .A(n2716), .ZN(n2682) );
  AOI222_X2 U1851 ( .A1(n3213), .A2(n460), .B1(n315), .B2(n457), .C1(n370), 
        .C2(n454), .ZN(n2716) );
  XOR2_X2 U1852 ( .A(n2683), .B(n265), .Z(n2036) );
  OAI21_X4 U1853 ( .B1(n2819), .B2(n339), .A(n2717), .ZN(n2683) );
  AOI222_X2 U1854 ( .A1(n3213), .A2(n457), .B1(n315), .B2(n454), .C1(n370), 
        .C2(n451), .ZN(n2717) );
  XOR2_X2 U1855 ( .A(n2684), .B(n265), .Z(n2037) );
  OAI21_X4 U1856 ( .B1(n2820), .B2(n339), .A(n2718), .ZN(n2684) );
  AOI222_X2 U1857 ( .A1(n3213), .A2(n454), .B1(n315), .B2(n451), .C1(n370), 
        .C2(n448), .ZN(n2718) );
  XOR2_X2 U1858 ( .A(n2685), .B(n265), .Z(n2038) );
  OAI21_X4 U1859 ( .B1(n2821), .B2(n339), .A(n2719), .ZN(n2685) );
  AOI222_X2 U1860 ( .A1(n3213), .A2(n451), .B1(n315), .B2(n448), .C1(n370), 
        .C2(n445), .ZN(n2719) );
  XOR2_X2 U1861 ( .A(n2686), .B(n265), .Z(n2039) );
  OAI21_X4 U1862 ( .B1(n2822), .B2(n339), .A(n2720), .ZN(n2686) );
  AOI222_X2 U1863 ( .A1(n3213), .A2(n448), .B1(n315), .B2(n445), .C1(n370), 
        .C2(n442), .ZN(n2720) );
  XOR2_X2 U1864 ( .A(n2687), .B(n265), .Z(n2040) );
  OAI21_X4 U1865 ( .B1(n2823), .B2(n339), .A(n2721), .ZN(n2687) );
  AOI222_X2 U1866 ( .A1(n3213), .A2(n445), .B1(n315), .B2(n442), .C1(n370), 
        .C2(n439), .ZN(n2721) );
  XOR2_X2 U1867 ( .A(n2688), .B(n265), .Z(n2041) );
  OAI21_X4 U1868 ( .B1(n2824), .B2(n339), .A(n2722), .ZN(n2688) );
  AOI222_X2 U1869 ( .A1(n3213), .A2(n442), .B1(n315), .B2(n439), .C1(n370), 
        .C2(n436), .ZN(n2722) );
  XOR2_X2 U1870 ( .A(n2689), .B(n265), .Z(n2042) );
  OAI21_X4 U1871 ( .B1(n2825), .B2(n339), .A(n2723), .ZN(n2689) );
  AOI222_X2 U1872 ( .A1(n3213), .A2(n439), .B1(n315), .B2(n436), .C1(n370), 
        .C2(n433), .ZN(n2723) );
  XOR2_X2 U1873 ( .A(n2690), .B(n265), .Z(n2043) );
  OAI21_X4 U1874 ( .B1(n2826), .B2(n339), .A(n2724), .ZN(n2690) );
  AOI222_X2 U1875 ( .A1(n3213), .A2(n436), .B1(n315), .B2(n433), .C1(n370), 
        .C2(n430), .ZN(n2724) );
  XOR2_X2 U1876 ( .A(n2691), .B(n265), .Z(n2044) );
  OAI21_X4 U1877 ( .B1(n2827), .B2(n339), .A(n2725), .ZN(n2691) );
  AOI222_X2 U1878 ( .A1(n3213), .A2(n433), .B1(n315), .B2(n430), .C1(n370), 
        .C2(n427), .ZN(n2725) );
  XOR2_X2 U1879 ( .A(n2692), .B(n265), .Z(n2045) );
  OAI21_X4 U1880 ( .B1(n2828), .B2(n339), .A(n2726), .ZN(n2692) );
  AOI222_X2 U1881 ( .A1(n3213), .A2(n430), .B1(n315), .B2(n427), .C1(n370), 
        .C2(n424), .ZN(n2726) );
  XOR2_X2 U1882 ( .A(n2693), .B(n265), .Z(n2046) );
  OAI21_X4 U1883 ( .B1(n2829), .B2(n339), .A(n2727), .ZN(n2693) );
  AOI222_X2 U1884 ( .A1(n3213), .A2(n427), .B1(n315), .B2(n424), .C1(n370), 
        .C2(n421), .ZN(n2727) );
  XOR2_X2 U1885 ( .A(n2694), .B(n265), .Z(n2047) );
  OAI21_X4 U1886 ( .B1(n2830), .B2(n339), .A(n2728), .ZN(n2694) );
  AOI222_X2 U1887 ( .A1(n3213), .A2(n424), .B1(n315), .B2(n421), .C1(n370), 
        .C2(n418), .ZN(n2728) );
  XOR2_X2 U1888 ( .A(n2695), .B(n265), .Z(n2048) );
  OAI21_X4 U1889 ( .B1(n2831), .B2(n339), .A(n2729), .ZN(n2695) );
  AOI222_X2 U1890 ( .A1(n3213), .A2(n421), .B1(n315), .B2(n418), .C1(n370), 
        .C2(n415), .ZN(n2729) );
  XOR2_X2 U1891 ( .A(n2696), .B(n265), .Z(n2049) );
  OAI21_X4 U1892 ( .B1(n2832), .B2(n339), .A(n2730), .ZN(n2696) );
  AOI222_X2 U1893 ( .A1(n3213), .A2(n418), .B1(n315), .B2(n415), .C1(n370), 
        .C2(n412), .ZN(n2730) );
  XOR2_X2 U1894 ( .A(n2697), .B(n265), .Z(n2050) );
  OAI21_X4 U1895 ( .B1(n2833), .B2(n339), .A(n2731), .ZN(n2697) );
  AOI222_X2 U1896 ( .A1(n3213), .A2(n415), .B1(n315), .B2(n412), .C1(n370), 
        .C2(n409), .ZN(n2731) );
  XOR2_X2 U1897 ( .A(n2698), .B(n265), .Z(n2051) );
  AOI222_X2 U1899 ( .A1(n3213), .A2(n412), .B1(n315), .B2(n409), .C1(n370), 
        .C2(n406), .ZN(n2732) );
  XOR2_X2 U1900 ( .A(n2699), .B(n265), .Z(n2052) );
  OAI21_X4 U1901 ( .B1(n2835), .B2(n339), .A(n2733), .ZN(n2699) );
  AOI222_X2 U1902 ( .A1(n3213), .A2(n409), .B1(n315), .B2(n406), .C1(n370), 
        .C2(n403), .ZN(n2733) );
  XOR2_X2 U1903 ( .A(n2700), .B(n265), .Z(n2053) );
  OAI21_X4 U1904 ( .B1(n2836), .B2(n339), .A(n2734), .ZN(n2700) );
  AOI222_X2 U1905 ( .A1(n3213), .A2(n406), .B1(n315), .B2(n403), .C1(n370), 
        .C2(n400), .ZN(n2734) );
  XOR2_X2 U1906 ( .A(n2701), .B(n265), .Z(n2054) );
  OAI21_X4 U1907 ( .B1(n2837), .B2(n339), .A(n2735), .ZN(n2701) );
  AOI222_X2 U1908 ( .A1(n3213), .A2(n403), .B1(n315), .B2(n400), .C1(n370), 
        .C2(n397), .ZN(n2735) );
  XOR2_X2 U1909 ( .A(n2702), .B(n265), .Z(n2055) );
  OAI21_X4 U1910 ( .B1(n2838), .B2(n339), .A(n2736), .ZN(n2702) );
  AOI222_X2 U1911 ( .A1(n3213), .A2(n400), .B1(n315), .B2(n397), .C1(n370), 
        .C2(n393), .ZN(n2736) );
  XOR2_X2 U1912 ( .A(n2703), .B(n265), .Z(n2056) );
  OAI21_X4 U1913 ( .B1(n2839), .B2(n339), .A(n2737), .ZN(n2703) );
  AOI222_X2 U1914 ( .A1(n3213), .A2(n397), .B1(n315), .B2(n393), .C1(n370), 
        .C2(n390), .ZN(n2737) );
  XOR2_X2 U1915 ( .A(n2704), .B(n265), .Z(n2057) );
  AND2_X4 U1921 ( .A1(n3213), .A2(n390), .ZN(n1403) );
  XOR2_X2 U1923 ( .A(n2740), .B(n262), .Z(n2060) );
  OAI21_X4 U1924 ( .B1(n2808), .B2(n336), .A(n2774), .ZN(n2740) );
  NAND2_X4 U1925 ( .A1(n368), .A2(n484), .ZN(n2774) );
  XOR2_X2 U1926 ( .A(n2741), .B(n262), .Z(n2061) );
  OAI21_X4 U1927 ( .B1(n2809), .B2(n336), .A(n2775), .ZN(n2741) );
  AOI21_X4 U1928 ( .B1(n368), .B2(n481), .A(n1404), .ZN(n2775) );
  AND2_X4 U1929 ( .A1(n313), .A2(n484), .ZN(n1404) );
  XOR2_X2 U1930 ( .A(n2742), .B(n262), .Z(n2062) );
  OAI21_X4 U1931 ( .B1(n2810), .B2(n336), .A(n2776), .ZN(n2742) );
  AOI222_X2 U1932 ( .A1(n3205), .A2(n484), .B1(n313), .B2(n481), .C1(n368), 
        .C2(n478), .ZN(n2776) );
  XOR2_X2 U1933 ( .A(n2743), .B(n262), .Z(n2063) );
  OAI21_X4 U1934 ( .B1(n2811), .B2(n336), .A(n2777), .ZN(n2743) );
  AOI222_X2 U1935 ( .A1(n3205), .A2(n481), .B1(n313), .B2(n478), .C1(n368), 
        .C2(n475), .ZN(n2777) );
  XOR2_X2 U1936 ( .A(n2744), .B(n262), .Z(n2064) );
  OAI21_X4 U1937 ( .B1(n2812), .B2(n336), .A(n2778), .ZN(n2744) );
  AOI222_X2 U1938 ( .A1(n3205), .A2(n478), .B1(n313), .B2(n475), .C1(n368), 
        .C2(n472), .ZN(n2778) );
  XOR2_X2 U1939 ( .A(n2745), .B(n262), .Z(n2065) );
  OAI21_X4 U1940 ( .B1(n2813), .B2(n336), .A(n2779), .ZN(n2745) );
  AOI222_X2 U1941 ( .A1(n3205), .A2(n475), .B1(n313), .B2(n472), .C1(n368), 
        .C2(n469), .ZN(n2779) );
  XOR2_X2 U1942 ( .A(n2746), .B(n262), .Z(n2066) );
  OAI21_X4 U1943 ( .B1(n2814), .B2(n336), .A(n2780), .ZN(n2746) );
  AOI222_X2 U1944 ( .A1(n3205), .A2(n472), .B1(n313), .B2(n469), .C1(n368), 
        .C2(n466), .ZN(n2780) );
  XOR2_X2 U1945 ( .A(n2747), .B(n262), .Z(n2067) );
  OAI21_X4 U1946 ( .B1(n2815), .B2(n336), .A(n2781), .ZN(n2747) );
  AOI222_X2 U1947 ( .A1(n3205), .A2(n469), .B1(n313), .B2(n466), .C1(n368), 
        .C2(n463), .ZN(n2781) );
  XOR2_X2 U1948 ( .A(n2748), .B(n262), .Z(n2068) );
  OAI21_X4 U1949 ( .B1(n2816), .B2(n336), .A(n2782), .ZN(n2748) );
  AOI222_X2 U1950 ( .A1(n3205), .A2(n466), .B1(n313), .B2(n463), .C1(n368), 
        .C2(n460), .ZN(n2782) );
  XOR2_X2 U1951 ( .A(n2749), .B(n262), .Z(n2069) );
  OAI21_X4 U1952 ( .B1(n2817), .B2(n336), .A(n2783), .ZN(n2749) );
  AOI222_X2 U1953 ( .A1(n3205), .A2(n463), .B1(n313), .B2(n460), .C1(n368), 
        .C2(n457), .ZN(n2783) );
  XOR2_X2 U1954 ( .A(n2750), .B(n262), .Z(n2070) );
  OAI21_X4 U1955 ( .B1(n2818), .B2(n336), .A(n2784), .ZN(n2750) );
  AOI222_X2 U1956 ( .A1(n3205), .A2(n460), .B1(n313), .B2(n457), .C1(n368), 
        .C2(n454), .ZN(n2784) );
  XOR2_X2 U1957 ( .A(n2751), .B(n262), .Z(n2071) );
  OAI21_X4 U1958 ( .B1(n2819), .B2(n336), .A(n2785), .ZN(n2751) );
  AOI222_X2 U1959 ( .A1(n3205), .A2(n457), .B1(n313), .B2(n454), .C1(n368), 
        .C2(n451), .ZN(n2785) );
  XOR2_X2 U1960 ( .A(n2752), .B(n262), .Z(n2072) );
  OAI21_X4 U1961 ( .B1(n2820), .B2(n336), .A(n2786), .ZN(n2752) );
  AOI222_X2 U1962 ( .A1(n3205), .A2(n454), .B1(n313), .B2(n451), .C1(n368), 
        .C2(n448), .ZN(n2786) );
  XOR2_X2 U1963 ( .A(n2753), .B(n262), .Z(n2073) );
  OAI21_X4 U1964 ( .B1(n2821), .B2(n336), .A(n2787), .ZN(n2753) );
  AOI222_X2 U1965 ( .A1(n3205), .A2(n451), .B1(n313), .B2(n448), .C1(n368), 
        .C2(n445), .ZN(n2787) );
  XOR2_X2 U1966 ( .A(n2754), .B(n262), .Z(n2074) );
  OAI21_X4 U1967 ( .B1(n2822), .B2(n336), .A(n2788), .ZN(n2754) );
  AOI222_X2 U1968 ( .A1(n3205), .A2(n448), .B1(n313), .B2(n445), .C1(n368), 
        .C2(n442), .ZN(n2788) );
  XOR2_X2 U1969 ( .A(n2755), .B(n262), .Z(n2075) );
  OAI21_X4 U1970 ( .B1(n2823), .B2(n336), .A(n2789), .ZN(n2755) );
  AOI222_X2 U1971 ( .A1(n3205), .A2(n445), .B1(n313), .B2(n442), .C1(n368), 
        .C2(n439), .ZN(n2789) );
  XOR2_X2 U1972 ( .A(n2756), .B(n262), .Z(n2076) );
  OAI21_X4 U1973 ( .B1(n2824), .B2(n336), .A(n2790), .ZN(n2756) );
  AOI222_X2 U1974 ( .A1(n3205), .A2(n442), .B1(n313), .B2(n439), .C1(n368), 
        .C2(n436), .ZN(n2790) );
  XOR2_X2 U1975 ( .A(n2757), .B(n262), .Z(n2077) );
  OAI21_X4 U1976 ( .B1(n2825), .B2(n336), .A(n2791), .ZN(n2757) );
  AOI222_X2 U1977 ( .A1(n3205), .A2(n439), .B1(n313), .B2(n436), .C1(n368), 
        .C2(n433), .ZN(n2791) );
  XOR2_X2 U1978 ( .A(n2758), .B(n262), .Z(n2078) );
  OAI21_X4 U1979 ( .B1(n2826), .B2(n336), .A(n2792), .ZN(n2758) );
  AOI222_X2 U1980 ( .A1(n3205), .A2(n436), .B1(n313), .B2(n433), .C1(n368), 
        .C2(n430), .ZN(n2792) );
  XOR2_X2 U1981 ( .A(n2759), .B(n262), .Z(n2079) );
  OAI21_X4 U1982 ( .B1(n2827), .B2(n336), .A(n2793), .ZN(n2759) );
  AOI222_X2 U1983 ( .A1(n3205), .A2(n433), .B1(n313), .B2(n430), .C1(n368), 
        .C2(n427), .ZN(n2793) );
  XOR2_X2 U1984 ( .A(n2760), .B(n262), .Z(n2080) );
  OAI21_X4 U1985 ( .B1(n2828), .B2(n336), .A(n2794), .ZN(n2760) );
  AOI222_X2 U1986 ( .A1(n3205), .A2(n430), .B1(n313), .B2(n427), .C1(n368), 
        .C2(n424), .ZN(n2794) );
  XOR2_X2 U1987 ( .A(n2761), .B(n262), .Z(n2081) );
  OAI21_X4 U1988 ( .B1(n2829), .B2(n336), .A(n2795), .ZN(n2761) );
  AOI222_X2 U1989 ( .A1(n3205), .A2(n427), .B1(n313), .B2(n424), .C1(n368), 
        .C2(n421), .ZN(n2795) );
  XOR2_X2 U1990 ( .A(n2762), .B(n262), .Z(n2082) );
  OAI21_X4 U1991 ( .B1(n2830), .B2(n336), .A(n2796), .ZN(n2762) );
  AOI222_X2 U1992 ( .A1(n3205), .A2(n424), .B1(n313), .B2(n421), .C1(n368), 
        .C2(n418), .ZN(n2796) );
  XOR2_X2 U1993 ( .A(n2763), .B(n262), .Z(n2083) );
  OAI21_X4 U1994 ( .B1(n2831), .B2(n336), .A(n2797), .ZN(n2763) );
  AOI222_X2 U1995 ( .A1(n3205), .A2(n421), .B1(n313), .B2(n418), .C1(n368), 
        .C2(n415), .ZN(n2797) );
  XOR2_X2 U1996 ( .A(n2764), .B(n262), .Z(n2084) );
  OAI21_X4 U1997 ( .B1(n2832), .B2(n336), .A(n2798), .ZN(n2764) );
  AOI222_X2 U1998 ( .A1(n3205), .A2(n418), .B1(n313), .B2(n415), .C1(n368), 
        .C2(n412), .ZN(n2798) );
  XOR2_X2 U1999 ( .A(n2765), .B(n262), .Z(n2085) );
  OAI21_X4 U2000 ( .B1(n2833), .B2(n336), .A(n2799), .ZN(n2765) );
  AOI222_X2 U2001 ( .A1(n3205), .A2(n415), .B1(n313), .B2(n412), .C1(n368), 
        .C2(n409), .ZN(n2799) );
  XOR2_X2 U2002 ( .A(n2766), .B(n262), .Z(n2086) );
  AOI222_X2 U2004 ( .A1(n3205), .A2(n412), .B1(n313), .B2(n409), .C1(n368), 
        .C2(n406), .ZN(n2800) );
  XOR2_X2 U2005 ( .A(n2767), .B(n262), .Z(n2087) );
  OAI21_X4 U2006 ( .B1(n2835), .B2(n336), .A(n2801), .ZN(n2767) );
  AOI222_X2 U2007 ( .A1(n3205), .A2(n409), .B1(n313), .B2(n406), .C1(n368), 
        .C2(n403), .ZN(n2801) );
  XOR2_X2 U2008 ( .A(n2768), .B(n262), .Z(n2088) );
  OAI21_X4 U2009 ( .B1(n2836), .B2(n336), .A(n2802), .ZN(n2768) );
  AOI222_X2 U2010 ( .A1(n3205), .A2(n406), .B1(n313), .B2(n403), .C1(n368), 
        .C2(n400), .ZN(n2802) );
  XOR2_X2 U2011 ( .A(n2769), .B(n262), .Z(n2089) );
  OAI21_X4 U2012 ( .B1(n2837), .B2(n336), .A(n2803), .ZN(n2769) );
  AOI222_X2 U2013 ( .A1(n3205), .A2(n403), .B1(n313), .B2(n400), .C1(n368), 
        .C2(n397), .ZN(n2803) );
  XOR2_X2 U2014 ( .A(n2770), .B(n262), .Z(n2090) );
  OAI21_X4 U2015 ( .B1(n2838), .B2(n336), .A(n2804), .ZN(n2770) );
  AOI222_X2 U2016 ( .A1(n3205), .A2(n400), .B1(n313), .B2(n397), .C1(n368), 
        .C2(n393), .ZN(n2804) );
  XOR2_X2 U2017 ( .A(n2771), .B(n262), .Z(n2091) );
  OAI21_X4 U2018 ( .B1(n2839), .B2(n336), .A(n2805), .ZN(n2771) );
  AOI222_X2 U2019 ( .A1(n3205), .A2(n397), .B1(n313), .B2(n393), .C1(n368), 
        .C2(n390), .ZN(n2805) );
  XOR2_X2 U2020 ( .A(n2772), .B(n262), .Z(n678) );
  OAI21_X4 U2021 ( .B1(n2840), .B2(n336), .A(n2806), .ZN(n2772) );
  OAI21_X4 U2024 ( .B1(n2841), .B2(n336), .A(n2807), .ZN(n2773) );
  AND2_X4 U2026 ( .A1(n3205), .A2(n390), .ZN(n1406) );
  AND3_X4 U2103 ( .A1(n2908), .A2(n2919), .A3(a[31]), .ZN(n388) );
  AND3_X4 U2107 ( .A1(n2931), .A2(n2909), .A3(n2920), .ZN(n386) );
  AND3_X4 U2112 ( .A1(n2932), .A2(n2910), .A3(n2921), .ZN(n384) );
  AND3_X4 U2117 ( .A1(n2933), .A2(n2911), .A3(n2922), .ZN(n382) );
  AND3_X4 U2122 ( .A1(n2934), .A2(n2912), .A3(n2923), .ZN(n380) );
  AND3_X4 U2127 ( .A1(n2935), .A2(n2913), .A3(n2924), .ZN(n378) );
  AND3_X4 U2132 ( .A1(n2936), .A2(n2914), .A3(n2925), .ZN(n376) );
  AND3_X4 U2137 ( .A1(n2937), .A2(n2915), .A3(n2926), .ZN(n374) );
  AND3_X4 U2152 ( .A1(n2940), .A2(n2929), .A3(n2918), .ZN(n368) );
  XNOR2_X2 U2158 ( .A(n1441), .B(n1440), .ZN(n2843) );
  NAND2_X4 U2159 ( .A1(n1441), .A2(n484), .ZN(n2808) );
  XOR2_X2 U2162 ( .A(n1452), .B(n1407), .Z(n2844) );
  OAI21_X4 U2163 ( .B1(n1600), .B2(n1442), .A(n1443), .ZN(n1441) );
  NAND2_X4 U2164 ( .A1(n1528), .A2(n1444), .ZN(n1442) );
  AOI21_X4 U2165 ( .B1(n1529), .B2(n1444), .A(n1445), .ZN(n1443) );
  NOR2_X4 U2166 ( .A1(n1488), .A2(n1446), .ZN(n1444) );
  OAI21_X4 U2167 ( .B1(n1489), .B2(n1446), .A(n1447), .ZN(n1445) );
  NAND2_X4 U2168 ( .A1(n1468), .A2(n1448), .ZN(n1446) );
  AOI21_X4 U2169 ( .B1(n1448), .B2(n1469), .A(n1449), .ZN(n1447) );
  NOR2_X4 U2170 ( .A1(n1459), .A2(n1450), .ZN(n1448) );
  OAI21_X4 U2171 ( .B1(n1450), .B2(n1462), .A(n1451), .ZN(n1449) );
  NAND2_X4 U2172 ( .A1(n1689), .A2(n1451), .ZN(n1407) );
  NOR2_X4 U2174 ( .A1(n481), .A2(n484), .ZN(n1450) );
  NAND2_X4 U2175 ( .A1(n481), .A2(n484), .ZN(n1451) );
  XOR2_X2 U2176 ( .A(n1463), .B(n1408), .Z(n2845) );
  AOI21_X4 U2177 ( .B1(n1599), .B2(n1453), .A(n1454), .ZN(n1452) );
  NOR2_X4 U2178 ( .A1(n1530), .A2(n1455), .ZN(n1453) );
  OAI21_X4 U2179 ( .B1(n1531), .B2(n1455), .A(n1456), .ZN(n1454) );
  NAND2_X4 U2180 ( .A1(n1457), .A2(n1490), .ZN(n1455) );
  AOI21_X4 U2181 ( .B1(n1457), .B2(n1491), .A(n1458), .ZN(n1456) );
  NOR2_X4 U2182 ( .A1(n1470), .A2(n1459), .ZN(n1457) );
  OAI21_X4 U2183 ( .B1(n1471), .B2(n1459), .A(n1462), .ZN(n1458) );
  NAND2_X4 U2186 ( .A1(n1690), .A2(n1462), .ZN(n1408) );
  NOR2_X4 U2188 ( .A1(n478), .A2(n481), .ZN(n1459) );
  NAND2_X4 U2189 ( .A1(n478), .A2(n481), .ZN(n1462) );
  XOR2_X2 U2190 ( .A(n1476), .B(n1409), .Z(n2846) );
  AOI21_X4 U2191 ( .B1(n1599), .B2(n1464), .A(n1465), .ZN(n1463) );
  NOR2_X4 U2192 ( .A1(n1530), .A2(n1466), .ZN(n1464) );
  OAI21_X4 U2193 ( .B1(n1531), .B2(n1466), .A(n1467), .ZN(n1465) );
  NAND2_X4 U2194 ( .A1(n1490), .A2(n1468), .ZN(n1466) );
  AOI21_X4 U2195 ( .B1(n1491), .B2(n1468), .A(n1469), .ZN(n1467) );
  NOR2_X4 U2200 ( .A1(n1483), .A2(n1474), .ZN(n1468) );
  OAI21_X4 U2201 ( .B1(n1474), .B2(n1484), .A(n1475), .ZN(n1469) );
  NAND2_X4 U2202 ( .A1(n1691), .A2(n1475), .ZN(n1409) );
  NOR2_X4 U2204 ( .A1(n475), .A2(n478), .ZN(n1474) );
  NAND2_X4 U2205 ( .A1(n475), .A2(n478), .ZN(n1475) );
  XOR2_X2 U2206 ( .A(n1485), .B(n1410), .Z(n2847) );
  AOI21_X4 U2207 ( .B1(n1599), .B2(n1477), .A(n1478), .ZN(n1476) );
  NOR2_X4 U2208 ( .A1(n1530), .A2(n1479), .ZN(n1477) );
  OAI21_X4 U2209 ( .B1(n1531), .B2(n1479), .A(n1480), .ZN(n1478) );
  NAND2_X4 U2210 ( .A1(n1490), .A2(n1692), .ZN(n1479) );
  AOI21_X4 U2211 ( .B1(n1491), .B2(n1692), .A(n1482), .ZN(n1480) );
  NAND2_X4 U2214 ( .A1(n1692), .A2(n1484), .ZN(n1410) );
  NOR2_X4 U2216 ( .A1(n472), .A2(n475), .ZN(n1483) );
  NAND2_X4 U2217 ( .A1(n472), .A2(n475), .ZN(n1484) );
  XOR2_X2 U2218 ( .A(n1498), .B(n1411), .Z(n2848) );
  AOI21_X4 U2219 ( .B1(n1599), .B2(n1486), .A(n1487), .ZN(n1485) );
  NOR2_X4 U2220 ( .A1(n1530), .A2(n1488), .ZN(n1486) );
  OAI21_X4 U2221 ( .B1(n1531), .B2(n1488), .A(n1489), .ZN(n1487) );
  NAND2_X4 U2226 ( .A1(n1512), .A2(n1494), .ZN(n1488) );
  AOI21_X4 U2227 ( .B1(n1494), .B2(n1513), .A(n1495), .ZN(n1489) );
  NOR2_X4 U2228 ( .A1(n1505), .A2(n1496), .ZN(n1494) );
  OAI21_X4 U2229 ( .B1(n1496), .B2(n1506), .A(n1497), .ZN(n1495) );
  NAND2_X4 U2230 ( .A1(n1693), .A2(n1497), .ZN(n1411) );
  NOR2_X4 U2232 ( .A1(n469), .A2(n472), .ZN(n1496) );
  NAND2_X4 U2233 ( .A1(n469), .A2(n472), .ZN(n1497) );
  XOR2_X2 U2234 ( .A(n1507), .B(n1412), .Z(n2849) );
  AOI21_X4 U2235 ( .B1(n1599), .B2(n1499), .A(n1500), .ZN(n1498) );
  NOR2_X4 U2236 ( .A1(n1530), .A2(n1501), .ZN(n1499) );
  OAI21_X4 U2237 ( .B1(n1531), .B2(n1501), .A(n1502), .ZN(n1500) );
  NAND2_X4 U2238 ( .A1(n1512), .A2(n1694), .ZN(n1501) );
  AOI21_X4 U2239 ( .B1(n1513), .B2(n1694), .A(n1504), .ZN(n1502) );
  NAND2_X4 U2242 ( .A1(n1694), .A2(n1506), .ZN(n1412) );
  NOR2_X4 U2244 ( .A1(n466), .A2(n469), .ZN(n1505) );
  NAND2_X4 U2245 ( .A1(n466), .A2(n469), .ZN(n1506) );
  XOR2_X2 U2246 ( .A(n1520), .B(n1413), .Z(n2850) );
  AOI21_X4 U2247 ( .B1(n1599), .B2(n1508), .A(n1509), .ZN(n1507) );
  NOR2_X4 U2248 ( .A1(n1530), .A2(n1510), .ZN(n1508) );
  OAI21_X4 U2249 ( .B1(n1531), .B2(n1510), .A(n1511), .ZN(n1509) );
  NOR2_X4 U2256 ( .A1(n1523), .A2(n1518), .ZN(n1512) );
  OAI21_X4 U2257 ( .B1(n1518), .B2(n1526), .A(n1519), .ZN(n1513) );
  NAND2_X4 U2258 ( .A1(n1695), .A2(n1519), .ZN(n1413) );
  NOR2_X4 U2260 ( .A1(n463), .A2(n466), .ZN(n1518) );
  NAND2_X4 U2261 ( .A1(n463), .A2(n466), .ZN(n1519) );
  XOR2_X2 U2262 ( .A(n1527), .B(n1414), .Z(n2851) );
  AOI21_X4 U2263 ( .B1(n1599), .B2(n1521), .A(n1522), .ZN(n1520) );
  NOR2_X4 U2264 ( .A1(n1530), .A2(n1523), .ZN(n1521) );
  OAI21_X4 U2265 ( .B1(n1531), .B2(n1523), .A(n1526), .ZN(n1522) );
  NAND2_X4 U2268 ( .A1(n1696), .A2(n1526), .ZN(n1414) );
  NOR2_X4 U2270 ( .A1(n460), .A2(n463), .ZN(n1523) );
  NAND2_X4 U2271 ( .A1(n460), .A2(n463), .ZN(n1526) );
  XOR2_X2 U2272 ( .A(n1540), .B(n1415), .Z(n2852) );
  AOI21_X4 U2273 ( .B1(n1599), .B2(n1528), .A(n1529), .ZN(n1527) );
  NOR2_X4 U2278 ( .A1(n1568), .A2(n1534), .ZN(n1528) );
  OAI21_X4 U2279 ( .B1(n1569), .B2(n1534), .A(n1535), .ZN(n1529) );
  NAND2_X4 U2280 ( .A1(n1552), .A2(n1536), .ZN(n1534) );
  AOI21_X4 U2281 ( .B1(n1536), .B2(n1555), .A(n1537), .ZN(n1535) );
  NOR2_X4 U2282 ( .A1(n1543), .A2(n1538), .ZN(n1536) );
  OAI21_X4 U2283 ( .B1(n1538), .B2(n1546), .A(n1539), .ZN(n1537) );
  NAND2_X4 U2284 ( .A1(n1697), .A2(n1539), .ZN(n1415) );
  NOR2_X4 U2286 ( .A1(n457), .A2(n460), .ZN(n1538) );
  NAND2_X4 U2287 ( .A1(n457), .A2(n460), .ZN(n1539) );
  XOR2_X2 U2288 ( .A(n1547), .B(n1416), .Z(n2853) );
  AOI21_X4 U2289 ( .B1(n1599), .B2(n1541), .A(n1542), .ZN(n1540) );
  NOR2_X4 U2290 ( .A1(n1550), .A2(n1543), .ZN(n1541) );
  OAI21_X4 U2291 ( .B1(n1551), .B2(n1543), .A(n1546), .ZN(n1542) );
  NAND2_X4 U2294 ( .A1(n1698), .A2(n1546), .ZN(n1416) );
  NOR2_X4 U2296 ( .A1(n454), .A2(n457), .ZN(n1543) );
  NAND2_X4 U2297 ( .A1(n454), .A2(n457), .ZN(n1546) );
  XOR2_X2 U2298 ( .A(n1558), .B(n1417), .Z(n2854) );
  AOI21_X4 U2299 ( .B1(n1599), .B2(n1548), .A(n1549), .ZN(n1547) );
  NAND2_X4 U2302 ( .A1(n1570), .A2(n1552), .ZN(n1550) );
  AOI21_X4 U2303 ( .B1(n1571), .B2(n1552), .A(n1555), .ZN(n1551) );
  NOR2_X4 U2306 ( .A1(n1561), .A2(n1556), .ZN(n1552) );
  OAI21_X4 U2307 ( .B1(n1556), .B2(n1564), .A(n1557), .ZN(n1555) );
  NAND2_X4 U2308 ( .A1(n1699), .A2(n1557), .ZN(n1417) );
  NOR2_X4 U2310 ( .A1(n451), .A2(n454), .ZN(n1556) );
  NAND2_X4 U2311 ( .A1(n451), .A2(n454), .ZN(n1557) );
  XOR2_X2 U2312 ( .A(n1565), .B(n1418), .Z(n2855) );
  AOI21_X4 U2313 ( .B1(n1599), .B2(n1559), .A(n1560), .ZN(n1558) );
  NOR2_X4 U2314 ( .A1(n1568), .A2(n1561), .ZN(n1559) );
  OAI21_X4 U2315 ( .B1(n1569), .B2(n1561), .A(n1564), .ZN(n1560) );
  NAND2_X4 U2318 ( .A1(n1700), .A2(n1564), .ZN(n1418) );
  NOR2_X4 U2320 ( .A1(n448), .A2(n451), .ZN(n1561) );
  NAND2_X4 U2321 ( .A1(n448), .A2(n451), .ZN(n1564) );
  XOR2_X2 U2322 ( .A(n1578), .B(n1419), .Z(n2856) );
  AOI21_X4 U2323 ( .B1(n1599), .B2(n1570), .A(n1571), .ZN(n1565) );
  NAND2_X4 U2330 ( .A1(n1586), .A2(n1574), .ZN(n1568) );
  AOI21_X4 U2331 ( .B1(n1574), .B2(n1587), .A(n1575), .ZN(n1569) );
  NOR2_X4 U2332 ( .A1(n1581), .A2(n1576), .ZN(n1574) );
  OAI21_X4 U2333 ( .B1(n1576), .B2(n1584), .A(n1577), .ZN(n1575) );
  NAND2_X4 U2334 ( .A1(n1701), .A2(n1577), .ZN(n1419) );
  NOR2_X4 U2336 ( .A1(n445), .A2(n448), .ZN(n1576) );
  NAND2_X4 U2337 ( .A1(n445), .A2(n448), .ZN(n1577) );
  XOR2_X2 U2338 ( .A(n1585), .B(n1420), .Z(n2857) );
  AOI21_X4 U2339 ( .B1(n1599), .B2(n1579), .A(n1580), .ZN(n1578) );
  NOR2_X4 U2340 ( .A1(n1588), .A2(n1581), .ZN(n1579) );
  OAI21_X4 U2341 ( .B1(n1589), .B2(n1581), .A(n1584), .ZN(n1580) );
  NAND2_X4 U2344 ( .A1(n1702), .A2(n1584), .ZN(n1420) );
  NOR2_X4 U2346 ( .A1(n442), .A2(n445), .ZN(n1581) );
  NAND2_X4 U2347 ( .A1(n442), .A2(n445), .ZN(n1584) );
  XOR2_X2 U2348 ( .A(n1594), .B(n1421), .Z(n2858) );
  AOI21_X4 U2349 ( .B1(n1599), .B2(n1586), .A(n1587), .ZN(n1585) );
  NOR2_X4 U2354 ( .A1(n1597), .A2(n1592), .ZN(n1586) );
  OAI21_X4 U2355 ( .B1(n1592), .B2(n1598), .A(n1593), .ZN(n1587) );
  NAND2_X4 U2356 ( .A1(n1703), .A2(n1593), .ZN(n1421) );
  NOR2_X4 U2358 ( .A1(n439), .A2(n442), .ZN(n1592) );
  NAND2_X4 U2359 ( .A1(n439), .A2(n442), .ZN(n1593) );
  XNOR2_X2 U2360 ( .A(n1599), .B(n1422), .ZN(n2859) );
  AOI21_X4 U2361 ( .B1(n1599), .B2(n1704), .A(n1596), .ZN(n1594) );
  NAND2_X4 U2364 ( .A1(n1704), .A2(n1598), .ZN(n1422) );
  NOR2_X4 U2366 ( .A1(n436), .A2(n439), .ZN(n1597) );
  NAND2_X4 U2367 ( .A1(n436), .A2(n439), .ZN(n1598) );
  XOR2_X2 U2368 ( .A(n1609), .B(n1423), .Z(n2860) );
  AOI21_X4 U2370 ( .B1(n1655), .B2(n1601), .A(n1602), .ZN(n1600) );
  NOR2_X4 U2371 ( .A1(n1629), .A2(n1603), .ZN(n1601) );
  OAI21_X4 U2372 ( .B1(n1630), .B2(n1603), .A(n1604), .ZN(n1602) );
  NAND2_X4 U2373 ( .A1(n1617), .A2(n1605), .ZN(n1603) );
  AOI21_X4 U2374 ( .B1(n1605), .B2(n1620), .A(n1606), .ZN(n1604) );
  NOR2_X4 U2375 ( .A1(n1612), .A2(n1607), .ZN(n1605) );
  OAI21_X4 U2376 ( .B1(n1607), .B2(n1613), .A(n1608), .ZN(n1606) );
  NAND2_X4 U2377 ( .A1(n1705), .A2(n1608), .ZN(n1423) );
  NOR2_X4 U2379 ( .A1(n433), .A2(n436), .ZN(n1607) );
  NAND2_X4 U2380 ( .A1(n433), .A2(n436), .ZN(n1608) );
  XNOR2_X2 U2381 ( .A(n1614), .B(n1424), .ZN(n2861) );
  AOI21_X4 U2382 ( .B1(n1614), .B2(n1706), .A(n1611), .ZN(n1609) );
  NAND2_X4 U2385 ( .A1(n1706), .A2(n1613), .ZN(n1424) );
  NOR2_X4 U2387 ( .A1(n430), .A2(n433), .ZN(n1612) );
  NAND2_X4 U2388 ( .A1(n430), .A2(n433), .ZN(n1613) );
  XOR2_X2 U2389 ( .A(n1623), .B(n1425), .Z(n2862) );
  OAI21_X4 U2390 ( .B1(n1654), .B2(n1615), .A(n1616), .ZN(n1614) );
  NAND2_X4 U2391 ( .A1(n1631), .A2(n1617), .ZN(n1615) );
  AOI21_X4 U2392 ( .B1(n1632), .B2(n1617), .A(n1620), .ZN(n1616) );
  NOR2_X4 U2395 ( .A1(n1626), .A2(n1621), .ZN(n1617) );
  OAI21_X4 U2396 ( .B1(n1621), .B2(n1627), .A(n1622), .ZN(n1620) );
  NAND2_X4 U2397 ( .A1(n1707), .A2(n1622), .ZN(n1425) );
  NOR2_X4 U2399 ( .A1(n427), .A2(n430), .ZN(n1621) );
  NAND2_X4 U2400 ( .A1(n427), .A2(n430), .ZN(n1622) );
  XNOR2_X2 U2401 ( .A(n1628), .B(n1426), .ZN(n2863) );
  AOI21_X4 U2402 ( .B1(n1628), .B2(n1708), .A(n1625), .ZN(n1623) );
  NAND2_X4 U2405 ( .A1(n1708), .A2(n1627), .ZN(n1426) );
  NOR2_X4 U2407 ( .A1(n424), .A2(n427), .ZN(n1626) );
  NAND2_X4 U2408 ( .A1(n424), .A2(n427), .ZN(n1627) );
  XOR2_X2 U2409 ( .A(n1639), .B(n1427), .Z(n2864) );
  OAI21_X4 U2410 ( .B1(n1654), .B2(n1629), .A(n1630), .ZN(n1628) );
  NAND2_X4 U2415 ( .A1(n1647), .A2(n1635), .ZN(n1629) );
  AOI21_X4 U2416 ( .B1(n1635), .B2(n1648), .A(n1636), .ZN(n1630) );
  NOR2_X4 U2417 ( .A1(n1642), .A2(n1637), .ZN(n1635) );
  OAI21_X4 U2418 ( .B1(n1637), .B2(n1643), .A(n1638), .ZN(n1636) );
  NAND2_X4 U2419 ( .A1(n1709), .A2(n1638), .ZN(n1427) );
  NOR2_X4 U2421 ( .A1(n421), .A2(n424), .ZN(n1637) );
  NAND2_X4 U2422 ( .A1(n421), .A2(n424), .ZN(n1638) );
  XNOR2_X2 U2423 ( .A(n1644), .B(n1428), .ZN(n2865) );
  AOI21_X4 U2424 ( .B1(n1644), .B2(n1710), .A(n1641), .ZN(n1639) );
  NAND2_X4 U2427 ( .A1(n1710), .A2(n1643), .ZN(n1428) );
  NOR2_X4 U2429 ( .A1(n418), .A2(n421), .ZN(n1642) );
  NAND2_X4 U2430 ( .A1(n418), .A2(n421), .ZN(n1643) );
  XNOR2_X2 U2431 ( .A(n1651), .B(n1429), .ZN(n2866) );
  OAI21_X4 U2432 ( .B1(n1654), .B2(n1645), .A(n1646), .ZN(n1644) );
  NOR2_X4 U2435 ( .A1(n1652), .A2(n1649), .ZN(n1647) );
  OAI21_X4 U2436 ( .B1(n1649), .B2(n1653), .A(n1650), .ZN(n1648) );
  NAND2_X4 U2437 ( .A1(n1711), .A2(n1650), .ZN(n1429) );
  NOR2_X4 U2439 ( .A1(n415), .A2(n418), .ZN(n1649) );
  NAND2_X4 U2440 ( .A1(n415), .A2(n418), .ZN(n1650) );
  XOR2_X2 U2441 ( .A(n1654), .B(n1430), .Z(n2867) );
  OAI21_X4 U2442 ( .B1(n1654), .B2(n1652), .A(n1653), .ZN(n1651) );
  NAND2_X4 U2443 ( .A1(n1712), .A2(n1653), .ZN(n1430) );
  NOR2_X4 U2445 ( .A1(n412), .A2(n415), .ZN(n1652) );
  NAND2_X4 U2446 ( .A1(n412), .A2(n415), .ZN(n1653) );
  XNOR2_X2 U2447 ( .A(n1662), .B(n1431), .ZN(n2868) );
  OAI21_X4 U2449 ( .B1(n1676), .B2(n1656), .A(n1657), .ZN(n1655) );
  NAND2_X4 U2450 ( .A1(n1666), .A2(n1658), .ZN(n1656) );
  AOI21_X4 U2451 ( .B1(n1658), .B2(n1667), .A(n1659), .ZN(n1657) );
  NOR2_X4 U2452 ( .A1(n1663), .A2(n1660), .ZN(n1658) );
  OAI21_X4 U2453 ( .B1(n1660), .B2(n1664), .A(n1661), .ZN(n1659) );
  NAND2_X4 U2454 ( .A1(n1713), .A2(n1661), .ZN(n1431) );
  NOR2_X4 U2456 ( .A1(n409), .A2(n412), .ZN(n1660) );
  NAND2_X4 U2457 ( .A1(n409), .A2(n412), .ZN(n1661) );
  XOR2_X2 U2458 ( .A(n1665), .B(n1432), .Z(n2869) );
  OAI21_X4 U2459 ( .B1(n1665), .B2(n1663), .A(n1664), .ZN(n1662) );
  NAND2_X4 U2460 ( .A1(n1714), .A2(n1664), .ZN(n1432) );
  NOR2_X4 U2462 ( .A1(n406), .A2(n409), .ZN(n1663) );
  NAND2_X4 U2463 ( .A1(n406), .A2(n409), .ZN(n1664) );
  XOR2_X2 U2464 ( .A(n1670), .B(n1433), .Z(n2870) );
  AOI21_X4 U2465 ( .B1(n1675), .B2(n1666), .A(n1667), .ZN(n1665) );
  NOR2_X4 U2466 ( .A1(n1673), .A2(n1668), .ZN(n1666) );
  OAI21_X4 U2467 ( .B1(n1668), .B2(n1674), .A(n1669), .ZN(n1667) );
  NAND2_X4 U2468 ( .A1(n1715), .A2(n1669), .ZN(n1433) );
  NOR2_X4 U2470 ( .A1(n403), .A2(n406), .ZN(n1668) );
  NAND2_X4 U2471 ( .A1(n403), .A2(n406), .ZN(n1669) );
  XNOR2_X2 U2472 ( .A(n1675), .B(n1434), .ZN(n2871) );
  AOI21_X4 U2473 ( .B1(n1675), .B2(n1716), .A(n1672), .ZN(n1670) );
  NAND2_X4 U2476 ( .A1(n1716), .A2(n1674), .ZN(n1434) );
  NOR2_X4 U2478 ( .A1(n400), .A2(n403), .ZN(n1673) );
  NAND2_X4 U2479 ( .A1(n400), .A2(n403), .ZN(n1674) );
  XNOR2_X2 U2480 ( .A(n1681), .B(n1435), .ZN(n2872) );
  AOI21_X4 U2482 ( .B1(n1677), .B2(n1685), .A(n1678), .ZN(n1676) );
  NOR2_X4 U2483 ( .A1(n1682), .A2(n1679), .ZN(n1677) );
  OAI21_X4 U2484 ( .B1(n1679), .B2(n1683), .A(n1680), .ZN(n1678) );
  NAND2_X4 U2485 ( .A1(n1717), .A2(n1680), .ZN(n1435) );
  NOR2_X4 U2487 ( .A1(n397), .A2(n400), .ZN(n1679) );
  NAND2_X4 U2488 ( .A1(n397), .A2(n400), .ZN(n1680) );
  XOR2_X2 U2489 ( .A(n1436), .B(n1684), .Z(n2873) );
  OAI21_X4 U2490 ( .B1(n1682), .B2(n1684), .A(n1683), .ZN(n1681) );
  NAND2_X4 U2491 ( .A1(n1718), .A2(n1683), .ZN(n1436) );
  NOR2_X4 U2493 ( .A1(n393), .A2(n397), .ZN(n1682) );
  NAND2_X4 U2494 ( .A1(n393), .A2(n397), .ZN(n1683) );
  NAND2_X4 U2498 ( .A1(n1719), .A2(n1684), .ZN(n2840) );
  NOR2_X4 U2500 ( .A1(n390), .A2(n393), .ZN(n1686) );
  NAND2_X4 U2501 ( .A1(n390), .A2(n393), .ZN(n1684) );
  INV_X1 U2506 ( .A(n268), .ZN(n3216) );
  INV_X1 U2507 ( .A(n271), .ZN(n3208) );
  INV_X1 U2508 ( .A(n262), .ZN(n3209) );
  XOR2_X1 U2509 ( .A(a[28]), .B(n289), .Z(n2931) );
  XNOR2_X1 U2510 ( .A(n277), .B(a[18]), .ZN(n2912) );
  XOR2_X1 U2511 ( .A(a[16]), .B(n277), .Z(n2935) );
  XNOR2_X1 U2512 ( .A(n286), .B(a[27]), .ZN(n2909) );
  XNOR2_X1 U2513 ( .A(a[27]), .B(a[28]), .ZN(n2920) );
  XOR2_X1 U2514 ( .A(a[25]), .B(n286), .Z(n2932) );
  XOR2_X1 U2515 ( .A(a[19]), .B(n280), .Z(n2934) );
  XNOR2_X1 U2516 ( .A(a[18]), .B(a[19]), .ZN(n2923) );
  XOR2_X1 U2517 ( .A(a[1]), .B(n262), .Z(n2940) );
  XNOR2_X1 U2518 ( .A(a[24]), .B(a[25]), .ZN(n2921) );
  XNOR2_X1 U2519 ( .A(n262), .B(a[3]), .ZN(n2917) );
  XOR2_X1 U2520 ( .A(a[4]), .B(n265), .Z(n2939) );
  XNOR2_X1 U2521 ( .A(a[3]), .B(a[4]), .ZN(n2928) );
  XOR2_X1 U2522 ( .A(a[22]), .B(n283), .Z(n2933) );
  XNOR2_X1 U2523 ( .A(a[21]), .B(a[22]), .ZN(n2922) );
  XNOR2_X1 U2524 ( .A(n265), .B(a[6]), .ZN(n2916) );
  XNOR2_X1 U2525 ( .A(a[6]), .B(a[7]), .ZN(n2927) );
  XNOR2_X1 U2526 ( .A(n271), .B(a[12]), .ZN(n2914) );
  XNOR2_X1 U2527 ( .A(n268), .B(a[9]), .ZN(n2915) );
  INV_X1 U2528 ( .A(a[10]), .ZN(n3210) );
  XNOR2_X1 U2529 ( .A(a[9]), .B(a[10]), .ZN(n2926) );
  XNOR2_X1 U2530 ( .A(n274), .B(a[15]), .ZN(n2913) );
  XNOR2_X1 U2531 ( .A(a[15]), .B(a[16]), .ZN(n2924) );
  XOR2_X1 U2532 ( .A(a[13]), .B(n274), .Z(n2936) );
  XNOR2_X1 U2533 ( .A(a[12]), .B(a[13]), .ZN(n2925) );
  XNOR2_X1 U2534 ( .A(a[0]), .B(a[1]), .ZN(n2929) );
  INV_X1 U2535 ( .A(a[0]), .ZN(n2918) );
  OR2_X1 U2536 ( .A1(n2929), .A2(a[0]), .ZN(n3227) );
  XNOR2_X1 U2537 ( .A(a[30]), .B(a[31]), .ZN(n2919) );
  AND3_X4 U2538 ( .A1(n2939), .A2(n2917), .A3(n2928), .ZN(n370) );
  OR2_X1 U2539 ( .A1(n2931), .A2(n2909), .ZN(n3126) );
  INV_X1 U2540 ( .A(n3126), .ZN(n3127) );
  INV_X1 U2541 ( .A(n3126), .ZN(n3128) );
  OR2_X1 U2542 ( .A1(n2908), .A2(a[31]), .ZN(n3129) );
  INV_X1 U2543 ( .A(n3129), .ZN(n3130) );
  INV_X1 U2544 ( .A(n3129), .ZN(n3131) );
  XNOR2_X1 U2545 ( .A(n289), .B(a[30]), .ZN(n2908) );
  OR2_X1 U2546 ( .A1(n2935), .A2(n2913), .ZN(n3132) );
  INV_X1 U2547 ( .A(n3132), .ZN(n3133) );
  INV_X1 U2548 ( .A(n3132), .ZN(n3134) );
  OR2_X1 U2549 ( .A1(n2934), .A2(n2912), .ZN(n3135) );
  INV_X1 U2550 ( .A(n3135), .ZN(n3136) );
  INV_X1 U2551 ( .A(n3135), .ZN(n3137) );
  OR2_X1 U2552 ( .A1(n2933), .A2(n2911), .ZN(n3138) );
  INV_X1 U2553 ( .A(n3138), .ZN(n3139) );
  INV_X1 U2554 ( .A(n3138), .ZN(n3140) );
  XNOR2_X1 U2555 ( .A(n280), .B(a[21]), .ZN(n2911) );
  NOR2_X4 U2556 ( .A1(n2932), .A2(n2910), .ZN(n3141) );
  XNOR2_X1 U2557 ( .A(n283), .B(a[24]), .ZN(n2910) );
  NOR2_X1 U2558 ( .A1(n2932), .A2(n2910), .ZN(n307) );
  NAND2_X4 U2559 ( .A1(n2931), .A2(n3218), .ZN(n363) );
  NAND2_X4 U2560 ( .A1(a[31]), .A2(n3217), .ZN(n366) );
  NAND2_X4 U2561 ( .A1(n2932), .A2(n3219), .ZN(n360) );
  XOR2_X1 U2562 ( .A(n773), .B(n782), .Z(n3142) );
  XOR2_X1 U2563 ( .A(n3142), .B(n531), .Z(product[51]) );
  NAND2_X1 U2564 ( .A1(n773), .A2(n782), .ZN(n3143) );
  NAND2_X1 U2565 ( .A1(n773), .A2(n531), .ZN(n3144) );
  NAND2_X1 U2566 ( .A1(n782), .A2(n531), .ZN(n3145) );
  NAND3_X1 U2567 ( .A1(n3143), .A2(n3144), .A3(n3145), .ZN(n530) );
  XOR2_X1 U2568 ( .A(n765), .B(n772), .Z(n3146) );
  XOR2_X1 U2569 ( .A(n3146), .B(n530), .Z(product[52]) );
  NAND2_X1 U2570 ( .A1(n765), .A2(n772), .ZN(n3147) );
  NAND2_X1 U2571 ( .A1(n765), .A2(n530), .ZN(n3148) );
  NAND2_X1 U2572 ( .A1(n772), .A2(n530), .ZN(n3149) );
  NAND3_X1 U2573 ( .A1(n3147), .A2(n3148), .A3(n3149), .ZN(n529) );
  XOR2_X1 U2574 ( .A(n926), .B(n943), .Z(n3150) );
  XOR2_X1 U2575 ( .A(n3150), .B(n543), .Z(product[39]) );
  NAND2_X2 U2576 ( .A1(n926), .A2(n943), .ZN(n3151) );
  NAND2_X1 U2577 ( .A1(n926), .A2(n543), .ZN(n3152) );
  NAND2_X1 U2578 ( .A1(n943), .A2(n543), .ZN(n3153) );
  NAND3_X2 U2579 ( .A1(n3151), .A2(n3152), .A3(n3153), .ZN(n542) );
  XOR2_X1 U2580 ( .A(n910), .B(n925), .Z(n3154) );
  XOR2_X1 U2581 ( .A(n3154), .B(n542), .Z(product[40]) );
  NAND2_X1 U2582 ( .A1(n910), .A2(n925), .ZN(n3155) );
  NAND2_X1 U2583 ( .A1(n910), .A2(n542), .ZN(n3156) );
  NAND2_X1 U2584 ( .A1(n925), .A2(n542), .ZN(n3157) );
  NAND3_X1 U2585 ( .A1(n3155), .A2(n3156), .A3(n3157), .ZN(n541) );
  AOI21_X1 U2586 ( .B1(n3161), .B2(n696), .A(n600), .ZN(n3158) );
  AOI21_X1 U2587 ( .B1(n595), .B2(n694), .A(n592), .ZN(n3159) );
  BUF_X1 U2588 ( .A(n643), .Z(n3160) );
  BUF_X1 U2589 ( .A(n603), .Z(n3161) );
  INV_X1 U2590 ( .A(n2938), .ZN(n3162) );
  INV_X1 U2591 ( .A(n3162), .ZN(n3163) );
  AOI21_X2 U2592 ( .B1(n603), .B2(n696), .A(n600), .ZN(n598) );
  OAI21_X1 U2593 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  AOI21_X2 U2594 ( .B1(n595), .B2(n694), .A(n592), .ZN(n590) );
  OAI21_X1 U2595 ( .B1(n644), .B2(n646), .A(n645), .ZN(n643) );
  OAI21_X1 U2596 ( .B1(n606), .B2(n604), .A(n605), .ZN(n603) );
  NOR2_X2 U2597 ( .A1(n1351), .A2(n1356), .ZN(n649) );
  AND2_X1 U2598 ( .A1(n2933), .A2(n3220), .ZN(n3164) );
  INV_X32 U2599 ( .A(n3164), .ZN(n357) );
  AND3_X1 U2600 ( .A1(n3163), .A2(n2916), .A3(n2927), .ZN(n372) );
  XOR2_X1 U2601 ( .A(n3158), .B(n498), .Z(product[22]) );
  XOR2_X1 U2602 ( .A(n630), .B(n506), .Z(product[14]) );
  XNOR2_X1 U2603 ( .A(n651), .B(n511), .ZN(product[9]) );
  XOR2_X1 U2604 ( .A(n614), .B(n502), .Z(product[18]) );
  OAI21_X1 U2605 ( .B1(n2834), .B2(n366), .A(n2120), .ZN(n1737) );
  OAI21_X1 U2606 ( .B1(n2834), .B2(n363), .A(n2188), .ZN(n2154) );
  OAI21_X1 U2607 ( .B1(n2834), .B2(n360), .A(n2256), .ZN(n2222) );
  OAI21_X1 U2608 ( .B1(n2834), .B2(n357), .A(n2324), .ZN(n2290) );
  OAI21_X1 U2609 ( .B1(n2834), .B2(n354), .A(n2392), .ZN(n2358) );
  OAI21_X1 U2610 ( .B1(n2834), .B2(n351), .A(n2460), .ZN(n2426) );
  OAI21_X1 U2611 ( .B1(n2834), .B2(n348), .A(n2528), .ZN(n2494) );
  OAI21_X1 U2612 ( .B1(n2834), .B2(n345), .A(n2596), .ZN(n2562) );
  OAI21_X1 U2613 ( .B1(n2834), .B2(n342), .A(n2664), .ZN(n2630) );
  OAI21_X1 U2614 ( .B1(n2834), .B2(n339), .A(n2732), .ZN(n2698) );
  OAI21_X1 U2615 ( .B1(n2834), .B2(n336), .A(n2800), .ZN(n2766) );
  AOI21_X4 U2616 ( .B1(n651), .B2(n708), .A(n648), .ZN(n646) );
  OAI21_X1 U2617 ( .B1(n2841), .B2(n339), .A(n2739), .ZN(n2705) );
  OAI21_X2 U2618 ( .B1(n558), .B2(n556), .A(n557), .ZN(n555) );
  XOR2_X1 U2619 ( .A(n558), .B(n488), .Z(product[32]) );
  XNOR2_X1 U2620 ( .A(n3161), .B(n499), .ZN(product[21]) );
  XOR2_X1 U2621 ( .A(n622), .B(n504), .Z(product[16]) );
  XNOR2_X1 U2622 ( .A(n635), .B(n507), .ZN(product[13]) );
  XOR2_X1 U2623 ( .A(n3159), .B(n496), .Z(product[24]) );
  INV_X2 U2624 ( .A(n299), .ZN(n3165) );
  INV_X8 U2625 ( .A(n3165), .ZN(n3166) );
  NOR2_X1 U2626 ( .A1(n2936), .A2(n2914), .ZN(n299) );
  INV_X1 U2627 ( .A(n633), .ZN(n704) );
  NAND3_X2 U2628 ( .A1(n3179), .A2(n3180), .A3(n3181), .ZN(n534) );
  OAI21_X2 U2629 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  INV_X2 U2630 ( .A(n372), .ZN(n3167) );
  INV_X1 U2631 ( .A(n3167), .ZN(n3168) );
  INV_X4 U2632 ( .A(n3167), .ZN(n3169) );
  XOR2_X1 U2633 ( .A(n582), .B(n494), .Z(product[26]) );
  NOR2_X1 U2634 ( .A1(n1323), .A2(n1330), .ZN(n633) );
  NAND2_X2 U2635 ( .A1(n1323), .A2(n1330), .ZN(n634) );
  XNOR2_X1 U2636 ( .A(n595), .B(n497), .ZN(product[23]) );
  NAND3_X2 U2637 ( .A1(n3171), .A2(n3172), .A3(n3173), .ZN(n524) );
  XOR2_X1 U2638 ( .A(n738), .B(n733), .Z(n3170) );
  XOR2_X1 U2639 ( .A(n3170), .B(n525), .Z(product[57]) );
  NAND2_X2 U2640 ( .A1(n738), .A2(n733), .ZN(n3171) );
  NAND2_X1 U2641 ( .A1(n738), .A2(n525), .ZN(n3172) );
  NAND2_X1 U2642 ( .A1(n733), .A2(n525), .ZN(n3173) );
  XOR2_X1 U2643 ( .A(n729), .B(n732), .Z(n3174) );
  XOR2_X1 U2644 ( .A(n3174), .B(n524), .Z(product[58]) );
  NAND2_X1 U2645 ( .A1(n729), .A2(n732), .ZN(n3175) );
  NAND2_X1 U2646 ( .A1(n729), .A2(n524), .ZN(n3176) );
  NAND2_X1 U2647 ( .A1(n732), .A2(n524), .ZN(n3177) );
  NAND3_X1 U2648 ( .A1(n3175), .A2(n3176), .A3(n3177), .ZN(n523) );
  XOR2_X1 U2649 ( .A(n814), .B(n824), .Z(n3178) );
  XOR2_X1 U2650 ( .A(n3178), .B(n535), .Z(product[47]) );
  NAND2_X2 U2651 ( .A1(n814), .A2(n824), .ZN(n3179) );
  NAND2_X1 U2652 ( .A1(n814), .A2(n535), .ZN(n3180) );
  NAND2_X1 U2653 ( .A1(n824), .A2(n535), .ZN(n3181) );
  XOR2_X1 U2654 ( .A(n802), .B(n813), .Z(n3182) );
  XOR2_X1 U2655 ( .A(n3182), .B(n534), .Z(product[48]) );
  NAND2_X1 U2656 ( .A1(n802), .A2(n813), .ZN(n3183) );
  NAND2_X1 U2657 ( .A1(n802), .A2(n534), .ZN(n3184) );
  NAND2_X1 U2658 ( .A1(n813), .A2(n534), .ZN(n3185) );
  NAND3_X1 U2659 ( .A1(n3183), .A2(n3184), .A3(n3185), .ZN(n533) );
  XOR2_X1 U2660 ( .A(n961), .B(n978), .Z(n3186) );
  XOR2_X1 U2661 ( .A(n3186), .B(n545), .Z(product[37]) );
  NAND2_X2 U2662 ( .A1(n961), .A2(n978), .ZN(n3187) );
  NAND2_X1 U2663 ( .A1(n961), .A2(n545), .ZN(n3188) );
  NAND2_X1 U2664 ( .A1(n978), .A2(n545), .ZN(n3189) );
  NAND3_X2 U2665 ( .A1(n3187), .A2(n3188), .A3(n3189), .ZN(n544) );
  XOR2_X1 U2666 ( .A(n944), .B(n960), .Z(n3190) );
  XOR2_X1 U2667 ( .A(n3190), .B(n544), .Z(product[38]) );
  NAND2_X1 U2668 ( .A1(n944), .A2(n960), .ZN(n3191) );
  NAND2_X1 U2669 ( .A1(n944), .A2(n544), .ZN(n3192) );
  NAND2_X1 U2670 ( .A1(n960), .A2(n544), .ZN(n3193) );
  NAND3_X1 U2671 ( .A1(n3191), .A2(n3192), .A3(n3193), .ZN(n543) );
  NAND2_X1 U2672 ( .A1(n519), .A2(n3214), .ZN(n3196) );
  NAND2_X1 U2673 ( .A1(n3194), .A2(n3195), .ZN(n3197) );
  NAND2_X1 U2674 ( .A1(n3196), .A2(n3197), .ZN(product[63]) );
  INV_X1 U2675 ( .A(n519), .ZN(n3194) );
  INV_X1 U2676 ( .A(n3214), .ZN(n3195) );
  BUF_X1 U2677 ( .A(n571), .Z(n3198) );
  BUF_X1 U2678 ( .A(n563), .Z(n3199) );
  BUF_X1 U2679 ( .A(n611), .Z(n3200) );
  BUF_X1 U2680 ( .A(n587), .Z(n3201) );
  BUF_X1 U2681 ( .A(n627), .Z(n3202) );
  BUF_X1 U2682 ( .A(n619), .Z(n3203) );
  INV_X1 U2683 ( .A(n485), .ZN(n3214) );
  INV_X2 U2684 ( .A(n291), .ZN(n3204) );
  INV_X8 U2685 ( .A(n3204), .ZN(n3205) );
  NOR2_X2 U2686 ( .A1(n2940), .A2(n2918), .ZN(n291) );
  INV_X1 U2687 ( .A(a[7]), .ZN(n3206) );
  OAI21_X2 U2688 ( .B1(n660), .B2(n662), .A(n661), .ZN(n659) );
  NAND2_X2 U2689 ( .A1(n2093), .A2(n262), .ZN(n682) );
  XNOR2_X2 U2690 ( .A(n3206), .B(n268), .ZN(n2938) );
  AND2_X4 U2691 ( .A1(n2939), .A2(n3226), .ZN(n3207) );
  INV_X32 U2692 ( .A(n3207), .ZN(n339) );
  OR2_X4 U2693 ( .A1(n2926), .A2(n3224), .ZN(n3230) );
  INV_X8 U2694 ( .A(n3230), .ZN(n319) );
  XNOR2_X1 U2695 ( .A(n2569), .B(n3208), .ZN(n1988) );
  XOR2_X1 U2696 ( .A(n2705), .B(n265), .Z(n2058) );
  NAND2_X4 U2697 ( .A1(n2934), .A2(n3221), .ZN(n354) );
  XNOR2_X2 U2698 ( .A(n2773), .B(n3209), .ZN(n2093) );
  OAI21_X1 U2699 ( .B1(n2841), .B2(n345), .A(n2603), .ZN(n2569) );
  AOI22_X1 U2700 ( .A1(n3213), .A2(n393), .B1(n315), .B2(n390), .ZN(n2738) );
  OAI21_X1 U2701 ( .B1(n2840), .B2(n339), .A(n2738), .ZN(n2704) );
  INV_X4 U2702 ( .A(n3228), .ZN(n315) );
  XNOR2_X2 U2703 ( .A(n3210), .B(n271), .ZN(n2937) );
  OR2_X4 U2704 ( .A1(n2937), .A2(n2915), .ZN(n3211) );
  INV_X32 U2705 ( .A(n3211), .ZN(n297) );
  AOI22_X1 U2706 ( .A1(n295), .A2(n393), .B1(n317), .B2(n390), .ZN(n2670) );
  OAI21_X1 U2707 ( .B1(n2840), .B2(n342), .A(n2670), .ZN(n2636) );
  INV_X8 U2708 ( .A(n3229), .ZN(n317) );
  NAND2_X4 U2709 ( .A1(n2935), .A2(n3222), .ZN(n351) );
  INV_X2 U2710 ( .A(n293), .ZN(n3212) );
  INV_X8 U2711 ( .A(n3212), .ZN(n3213) );
  NOR2_X1 U2712 ( .A1(n2939), .A2(n2917), .ZN(n293) );
  OR2_X4 U2713 ( .A1(n2938), .A2(n2916), .ZN(n3215) );
  INV_X32 U2714 ( .A(n3215), .ZN(n295) );
  XNOR2_X1 U2715 ( .A(n2637), .B(n3216), .ZN(n2023) );
  AOI21_X4 U2716 ( .B1(n579), .B2(n690), .A(n576), .ZN(n574) );
  AOI21_X4 U2717 ( .B1(n571), .B2(n688), .A(n568), .ZN(n566) );
  XNOR2_X1 U2718 ( .A(n3199), .B(n489), .ZN(product[31]) );
  XNOR2_X1 U2719 ( .A(n3200), .B(n501), .ZN(product[19]) );
  XNOR2_X1 U2720 ( .A(n3203), .B(n503), .ZN(product[17]) );
  XOR2_X1 U2721 ( .A(n566), .B(n490), .Z(product[30]) );
  OAI21_X2 U2722 ( .B1(n566), .B2(n564), .A(n565), .ZN(n563) );
  NAND2_X4 U2723 ( .A1(n2936), .A2(n3223), .ZN(n348) );
  OAI21_X2 U2724 ( .B1(n614), .B2(n612), .A(n613), .ZN(n611) );
  NAND2_X4 U2725 ( .A1(n2940), .A2(a[0]), .ZN(n336) );
  OAI21_X2 U2726 ( .B1(n622), .B2(n620), .A(n621), .ZN(n619) );
  NAND2_X4 U2727 ( .A1(n2937), .A2(n3224), .ZN(n345) );
  XNOR2_X1 U2728 ( .A(n3160), .B(n509), .ZN(product[11]) );
  XNOR2_X1 U2729 ( .A(n3198), .B(n491), .ZN(product[29]) );
  XOR2_X1 U2730 ( .A(n550), .B(n486), .Z(product[34]) );
  XNOR2_X1 U2731 ( .A(n579), .B(n493), .ZN(product[27]) );
  XNOR2_X1 U2732 ( .A(n3202), .B(n505), .ZN(product[15]) );
  XNOR2_X1 U2733 ( .A(n555), .B(n487), .ZN(product[33]) );
  XNOR2_X1 U2734 ( .A(n3201), .B(n495), .ZN(product[25]) );
  XOR2_X1 U2735 ( .A(n574), .B(n492), .Z(product[28]) );
  XOR2_X1 U2736 ( .A(n510), .B(n646), .Z(product[10]) );
  AOI21_X2 U2737 ( .B1(n555), .B2(n684), .A(n552), .ZN(n550) );
  OAI21_X2 U2738 ( .B1(n574), .B2(n572), .A(n573), .ZN(n571) );
  OAI21_X1 U2739 ( .B1(n2841), .B2(n342), .A(n2671), .ZN(n2637) );
  NAND2_X4 U2740 ( .A1(n3163), .A2(n3225), .ZN(n342) );
  OAI21_X1 U2741 ( .B1(n550), .B2(n548), .A(n549), .ZN(n547) );
  OAI21_X2 U2742 ( .B1(n582), .B2(n580), .A(n581), .ZN(n579) );
  OAI21_X2 U2743 ( .B1(n590), .B2(n588), .A(n589), .ZN(n587) );
  OAI21_X2 U2744 ( .B1(n630), .B2(n628), .A(n629), .ZN(n627) );
  OAI21_X2 U2745 ( .B1(n654), .B2(n652), .A(n653), .ZN(n651) );
  INV_X2 U2746 ( .A(n518), .ZN(product[0]) );
  INV_X2 U2747 ( .A(n941), .ZN(n959) );
  INV_X2 U2748 ( .A(n907), .ZN(n908) );
  INV_X2 U2749 ( .A(n891), .ZN(n892) );
  INV_X2 U2750 ( .A(n848), .ZN(n862) );
  INV_X2 U2751 ( .A(n811), .ZN(n823) );
  INV_X2 U2752 ( .A(n780), .ZN(n790) );
  INV_X2 U2753 ( .A(n755), .ZN(n763) );
  INV_X2 U2754 ( .A(n736), .ZN(n742) );
  INV_X2 U2755 ( .A(n723), .ZN(n727) );
  INV_X2 U2756 ( .A(n717), .ZN(n718) );
  INV_X2 U2757 ( .A(n1720), .ZN(n716) );
  INV_X2 U2758 ( .A(n681), .ZN(n715) );
  INV_X2 U2759 ( .A(n668), .ZN(n713) );
  INV_X2 U2760 ( .A(n660), .ZN(n711) );
  INV_X2 U2761 ( .A(n652), .ZN(n709) );
  INV_X2 U2762 ( .A(n644), .ZN(n707) );
  INV_X2 U2763 ( .A(n636), .ZN(n705) );
  INV_X2 U2764 ( .A(n628), .ZN(n703) );
  INV_X2 U2765 ( .A(n620), .ZN(n701) );
  INV_X2 U2766 ( .A(n612), .ZN(n699) );
  INV_X2 U2767 ( .A(n604), .ZN(n697) );
  INV_X2 U2768 ( .A(n596), .ZN(n695) );
  INV_X2 U2769 ( .A(n588), .ZN(n693) );
  INV_X2 U2770 ( .A(n580), .ZN(n691) );
  INV_X2 U2771 ( .A(n572), .ZN(n689) );
  INV_X2 U2772 ( .A(n564), .ZN(n687) );
  INV_X2 U2773 ( .A(n556), .ZN(n685) );
  INV_X2 U2774 ( .A(n548), .ZN(n683) );
  INV_X2 U2775 ( .A(n682), .ZN(n680) );
  INV_X2 U2776 ( .A(n678), .ZN(n679) );
  INV_X2 U2777 ( .A(n2091), .ZN(n676) );
  INV_X2 U2778 ( .A(n674), .ZN(n672) );
  INV_X2 U2779 ( .A(n673), .ZN(n714) );
  INV_X2 U2780 ( .A(n666), .ZN(n664) );
  INV_X2 U2781 ( .A(n665), .ZN(n712) );
  INV_X2 U2782 ( .A(n658), .ZN(n656) );
  INV_X2 U2783 ( .A(n657), .ZN(n710) );
  INV_X2 U2784 ( .A(n650), .ZN(n648) );
  INV_X2 U2785 ( .A(n649), .ZN(n708) );
  INV_X2 U2786 ( .A(n642), .ZN(n640) );
  INV_X2 U2787 ( .A(n641), .ZN(n706) );
  INV_X2 U2788 ( .A(n634), .ZN(n632) );
  INV_X2 U2789 ( .A(n626), .ZN(n624) );
  INV_X2 U2790 ( .A(n625), .ZN(n702) );
  INV_X2 U2791 ( .A(n618), .ZN(n616) );
  INV_X2 U2792 ( .A(n617), .ZN(n700) );
  INV_X2 U2793 ( .A(n610), .ZN(n608) );
  INV_X2 U2794 ( .A(n609), .ZN(n698) );
  INV_X2 U2795 ( .A(n602), .ZN(n600) );
  INV_X2 U2796 ( .A(n601), .ZN(n696) );
  INV_X2 U2797 ( .A(n594), .ZN(n592) );
  INV_X2 U2798 ( .A(n593), .ZN(n694) );
  INV_X2 U2799 ( .A(n586), .ZN(n584) );
  INV_X2 U2800 ( .A(n585), .ZN(n692) );
  INV_X2 U2801 ( .A(n578), .ZN(n576) );
  INV_X2 U2802 ( .A(n577), .ZN(n690) );
  INV_X2 U2803 ( .A(n570), .ZN(n568) );
  INV_X2 U2804 ( .A(n569), .ZN(n688) );
  INV_X2 U2805 ( .A(n562), .ZN(n560) );
  INV_X2 U2806 ( .A(n561), .ZN(n686) );
  INV_X2 U2807 ( .A(n554), .ZN(n552) );
  INV_X2 U2808 ( .A(n553), .ZN(n684) );
  INV_X2 U2809 ( .A(n390), .ZN(n2841) );
  INV_X2 U2810 ( .A(n2873), .ZN(n2839) );
  INV_X2 U2811 ( .A(n2872), .ZN(n2838) );
  INV_X2 U2812 ( .A(n2871), .ZN(n2837) );
  INV_X2 U2813 ( .A(n2870), .ZN(n2836) );
  INV_X2 U2814 ( .A(n2869), .ZN(n2835) );
  INV_X2 U2815 ( .A(n2868), .ZN(n2834) );
  INV_X2 U2816 ( .A(n2867), .ZN(n2833) );
  INV_X2 U2817 ( .A(n2866), .ZN(n2832) );
  INV_X2 U2818 ( .A(n2865), .ZN(n2831) );
  INV_X2 U2819 ( .A(n2864), .ZN(n2830) );
  INV_X2 U2820 ( .A(n2863), .ZN(n2829) );
  INV_X2 U2821 ( .A(n2862), .ZN(n2828) );
  INV_X2 U2822 ( .A(n2861), .ZN(n2827) );
  INV_X2 U2823 ( .A(n2860), .ZN(n2826) );
  INV_X2 U2824 ( .A(n2859), .ZN(n2825) );
  INV_X2 U2825 ( .A(n2858), .ZN(n2824) );
  INV_X2 U2826 ( .A(n2857), .ZN(n2823) );
  INV_X2 U2827 ( .A(n2856), .ZN(n2822) );
  INV_X2 U2828 ( .A(n2855), .ZN(n2821) );
  INV_X2 U2829 ( .A(n2854), .ZN(n2820) );
  INV_X2 U2830 ( .A(n2853), .ZN(n2819) );
  INV_X2 U2831 ( .A(n2852), .ZN(n2818) );
  INV_X2 U2832 ( .A(n2851), .ZN(n2817) );
  INV_X2 U2833 ( .A(n2850), .ZN(n2816) );
  INV_X2 U2834 ( .A(n2849), .ZN(n2815) );
  INV_X2 U2835 ( .A(n2848), .ZN(n2814) );
  INV_X2 U2836 ( .A(n2847), .ZN(n2813) );
  INV_X2 U2837 ( .A(n2846), .ZN(n2812) );
  INV_X2 U2838 ( .A(n2845), .ZN(n2811) );
  INV_X2 U2839 ( .A(n2844), .ZN(n2810) );
  INV_X2 U2840 ( .A(n2843), .ZN(n2809) );
  INV_X2 U2841 ( .A(n1406), .ZN(n2807) );
  AOI22_X2 U2842 ( .A1(n3205), .A2(n393), .B1(n313), .B2(n390), .ZN(n2806) );
  INV_X2 U2843 ( .A(n3227), .ZN(n313) );
  INV_X2 U2844 ( .A(n1403), .ZN(n2739) );
  OR2_X2 U2845 ( .A1(n2928), .A2(n3226), .ZN(n3228) );
  INV_X2 U2846 ( .A(n2917), .ZN(n3226) );
  INV_X2 U2847 ( .A(n1400), .ZN(n2671) );
  OR2_X2 U2848 ( .A1(n2927), .A2(n3225), .ZN(n3229) );
  INV_X2 U2849 ( .A(n2916), .ZN(n3225) );
  INV_X2 U2850 ( .A(n1397), .ZN(n2603) );
  AOI22_X2 U2851 ( .A1(n297), .A2(n393), .B1(n319), .B2(n390), .ZN(n2602) );
  INV_X2 U2852 ( .A(n2915), .ZN(n3224) );
  INV_X2 U2853 ( .A(n1394), .ZN(n2535) );
  AOI22_X2 U2854 ( .A1(n3166), .A2(n393), .B1(n321), .B2(n390), .ZN(n2534) );
  INV_X2 U2855 ( .A(n3231), .ZN(n321) );
  OR2_X2 U2856 ( .A1(n2925), .A2(n3223), .ZN(n3231) );
  INV_X2 U2857 ( .A(n2914), .ZN(n3223) );
  INV_X2 U2858 ( .A(n1391), .ZN(n2467) );
  AOI22_X2 U2859 ( .A1(n3134), .A2(n393), .B1(n323), .B2(n390), .ZN(n2466) );
  INV_X2 U2860 ( .A(n3232), .ZN(n323) );
  OR2_X2 U2861 ( .A1(n2924), .A2(n3222), .ZN(n3232) );
  INV_X2 U2862 ( .A(n2913), .ZN(n3222) );
  INV_X2 U2863 ( .A(n1388), .ZN(n2399) );
  AOI22_X2 U2864 ( .A1(n3137), .A2(n393), .B1(n325), .B2(n390), .ZN(n2398) );
  INV_X2 U2865 ( .A(n3233), .ZN(n325) );
  OR2_X2 U2866 ( .A1(n2923), .A2(n3221), .ZN(n3233) );
  INV_X2 U2867 ( .A(n2912), .ZN(n3221) );
  INV_X2 U2868 ( .A(n1385), .ZN(n2331) );
  AOI22_X2 U2869 ( .A1(n3140), .A2(n393), .B1(n327), .B2(n390), .ZN(n2330) );
  INV_X2 U2870 ( .A(n3234), .ZN(n327) );
  OR2_X2 U2871 ( .A1(n2922), .A2(n3220), .ZN(n3234) );
  INV_X2 U2872 ( .A(n2911), .ZN(n3220) );
  INV_X2 U2873 ( .A(n1382), .ZN(n2263) );
  AOI22_X2 U2874 ( .A1(n307), .A2(n393), .B1(n329), .B2(n390), .ZN(n2262) );
  INV_X2 U2875 ( .A(n3235), .ZN(n329) );
  OR2_X2 U2876 ( .A1(n2921), .A2(n3219), .ZN(n3235) );
  INV_X2 U2877 ( .A(n2910), .ZN(n3219) );
  INV_X2 U2878 ( .A(n1379), .ZN(n2195) );
  AOI22_X2 U2879 ( .A1(n3128), .A2(n393), .B1(n331), .B2(n390), .ZN(n2194) );
  INV_X2 U2880 ( .A(n3236), .ZN(n331) );
  OR2_X2 U2881 ( .A1(n2920), .A2(n3218), .ZN(n3236) );
  INV_X2 U2882 ( .A(n2909), .ZN(n3218) );
  INV_X2 U2883 ( .A(n1376), .ZN(n2127) );
  AOI22_X2 U2884 ( .A1(n3130), .A2(n393), .B1(n333), .B2(n390), .ZN(n2126) );
  INV_X2 U2885 ( .A(n3237), .ZN(n333) );
  OR2_X2 U2886 ( .A1(n2919), .A2(n3217), .ZN(n3237) );
  INV_X2 U2887 ( .A(n2908), .ZN(n3217) );
  INV_X2 U2888 ( .A(n265), .ZN(n2024) );
  INV_X2 U2889 ( .A(n274), .ZN(n1919) );
  INV_X2 U2890 ( .A(n277), .ZN(n1884) );
  INV_X2 U2891 ( .A(n280), .ZN(n1849) );
  INV_X2 U2892 ( .A(n283), .ZN(n1814) );
  INV_X2 U2893 ( .A(n286), .ZN(n1779) );
  INV_X2 U2894 ( .A(n289), .ZN(n1745) );
  INV_X2 U2895 ( .A(n1686), .ZN(n1719) );
  INV_X2 U2896 ( .A(n1682), .ZN(n1718) );
  INV_X2 U2897 ( .A(n1679), .ZN(n1717) );
  INV_X2 U2898 ( .A(n1668), .ZN(n1715) );
  INV_X2 U2899 ( .A(n1663), .ZN(n1714) );
  INV_X2 U2900 ( .A(n1660), .ZN(n1713) );
  INV_X2 U2901 ( .A(n1652), .ZN(n1712) );
  INV_X2 U2902 ( .A(n1649), .ZN(n1711) );
  INV_X2 U2903 ( .A(n1637), .ZN(n1709) );
  INV_X2 U2904 ( .A(n1621), .ZN(n1707) );
  INV_X2 U2905 ( .A(n1607), .ZN(n1705) );
  INV_X2 U2906 ( .A(n1592), .ZN(n1703) );
  INV_X2 U2907 ( .A(n1581), .ZN(n1702) );
  INV_X2 U2908 ( .A(n1576), .ZN(n1701) );
  INV_X2 U2909 ( .A(n1561), .ZN(n1700) );
  INV_X2 U2910 ( .A(n1556), .ZN(n1699) );
  INV_X2 U2911 ( .A(n1543), .ZN(n1698) );
  INV_X2 U2912 ( .A(n1538), .ZN(n1697) );
  INV_X2 U2913 ( .A(n1523), .ZN(n1696) );
  INV_X2 U2914 ( .A(n1518), .ZN(n1695) );
  INV_X2 U2915 ( .A(n1496), .ZN(n1693) );
  INV_X2 U2916 ( .A(n1474), .ZN(n1691) );
  INV_X2 U2917 ( .A(n1459), .ZN(n1690) );
  INV_X2 U2918 ( .A(n1450), .ZN(n1689) );
  INV_X2 U2919 ( .A(n1684), .ZN(n1685) );
  INV_X2 U2920 ( .A(n1676), .ZN(n1675) );
  INV_X2 U2921 ( .A(n1674), .ZN(n1672) );
  INV_X2 U2922 ( .A(n1673), .ZN(n1716) );
  INV_X2 U2923 ( .A(n1655), .ZN(n1654) );
  INV_X2 U2924 ( .A(n1648), .ZN(n1646) );
  INV_X2 U2925 ( .A(n1647), .ZN(n1645) );
  INV_X2 U2926 ( .A(n1643), .ZN(n1641) );
  INV_X2 U2927 ( .A(n1642), .ZN(n1710) );
  INV_X2 U2928 ( .A(n1630), .ZN(n1632) );
  INV_X2 U2929 ( .A(n1629), .ZN(n1631) );
  INV_X2 U2930 ( .A(n1627), .ZN(n1625) );
  INV_X2 U2931 ( .A(n1626), .ZN(n1708) );
  INV_X2 U2932 ( .A(n1613), .ZN(n1611) );
  INV_X2 U2933 ( .A(n1612), .ZN(n1706) );
  INV_X2 U2934 ( .A(n1600), .ZN(n1599) );
  INV_X2 U2935 ( .A(n1598), .ZN(n1596) );
  INV_X2 U2936 ( .A(n1597), .ZN(n1704) );
  INV_X2 U2937 ( .A(n1587), .ZN(n1589) );
  INV_X2 U2938 ( .A(n1586), .ZN(n1588) );
  INV_X2 U2939 ( .A(n1569), .ZN(n1571) );
  INV_X2 U2940 ( .A(n1568), .ZN(n1570) );
  INV_X2 U2941 ( .A(n1551), .ZN(n1549) );
  INV_X2 U2942 ( .A(n1550), .ZN(n1548) );
  INV_X2 U2943 ( .A(n1529), .ZN(n1531) );
  INV_X2 U2944 ( .A(n1528), .ZN(n1530) );
  INV_X2 U2945 ( .A(n1513), .ZN(n1511) );
  INV_X2 U2946 ( .A(n1512), .ZN(n1510) );
  INV_X2 U2947 ( .A(n1506), .ZN(n1504) );
  INV_X2 U2948 ( .A(n1505), .ZN(n1694) );
  INV_X2 U2949 ( .A(n1489), .ZN(n1491) );
  INV_X2 U2950 ( .A(n1488), .ZN(n1490) );
  INV_X2 U2951 ( .A(n1484), .ZN(n1482) );
  INV_X2 U2952 ( .A(n1483), .ZN(n1692) );
  INV_X2 U2953 ( .A(n1469), .ZN(n1471) );
  INV_X2 U2954 ( .A(n1468), .ZN(n1470) );
  INV_X2 U2955 ( .A(n484), .ZN(n1440) );
endmodule


module mul32_0_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n262, n265, n268, n271, n274, n277, n280, n283, n286, n289, n291,
         n293, n295, n297, n303, n313, n315, n317, n319, n321, n323, n325,
         n327, n329, n331, n333, n336, n339, n342, n345, n348, n351, n354,
         n357, n368, n370, n372, n374, n376, n378, n380, n382, n384, n386,
         n388, n390, n393, n397, n400, n403, n406, n409, n412, n415, n418,
         n421, n424, n427, n430, n433, n436, n439, n442, n445, n448, n451,
         n454, n457, n460, n463, n466, n469, n472, n475, n478, n481, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n552, n553, n554, n555, n556, n557, n558, n560, n561, n562, n563,
         n564, n565, n566, n568, n569, n570, n571, n572, n573, n574, n576,
         n577, n578, n579, n580, n581, n582, n584, n585, n586, n587, n588,
         n589, n590, n592, n593, n594, n595, n596, n597, n598, n600, n601,
         n602, n603, n604, n605, n606, n608, n609, n610, n611, n612, n613,
         n614, n616, n617, n618, n619, n620, n621, n622, n624, n625, n626,
         n627, n628, n629, n630, n632, n633, n634, n635, n636, n637, n638,
         n640, n641, n642, n643, n644, n645, n646, n648, n649, n650, n651,
         n652, n653, n654, n656, n657, n658, n659, n660, n661, n662, n664,
         n665, n666, n667, n668, n669, n670, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1376, n1377, n1379, n1380, n1382, n1383, n1385, n1386,
         n1388, n1389, n1391, n1392, n1394, n1395, n1397, n1398, n1400, n1401,
         n1403, n1404, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1518,
         n1519, n1520, n1521, n1522, n1523, n1526, n1527, n1528, n1529, n1530,
         n1531, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1564, n1565, n1568, n1569, n1570,
         n1571, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1584,
         n1585, n1586, n1587, n1588, n1589, n1592, n1593, n1594, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1620,
         n1621, n1622, n1623, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1635, n1636, n1637, n1638, n1639, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255;
  assign n262 = a[2];
  assign n265 = a[5];
  assign n268 = a[8];
  assign n271 = a[11];
  assign n274 = a[14];
  assign n277 = a[17];
  assign n280 = a[20];
  assign n283 = a[23];
  assign n286 = a[26];
  assign n289 = a[29];
  assign n390 = b[0];
  assign n393 = b[1];
  assign n397 = b[2];
  assign n400 = b[3];
  assign n403 = b[4];
  assign n406 = b[5];
  assign n409 = b[6];
  assign n412 = b[7];
  assign n415 = b[8];
  assign n418 = b[9];
  assign n421 = b[10];
  assign n424 = b[11];
  assign n427 = b[12];
  assign n430 = b[13];
  assign n433 = b[14];
  assign n436 = b[15];
  assign n439 = b[16];
  assign n442 = b[17];
  assign n445 = b[18];
  assign n448 = b[19];
  assign n451 = b[20];
  assign n454 = b[21];
  assign n457 = b[22];
  assign n460 = b[23];
  assign n463 = b[24];
  assign n466 = b[25];
  assign n469 = b[26];
  assign n472 = b[27];
  assign n475 = b[28];
  assign n478 = b[29];
  assign n481 = b[30];
  assign n484 = b[31];

  XOR2_X2 U304 ( .A(n717), .B(n716), .Z(n485) );
  FA_X1 U306 ( .A(n720), .B(n721), .CI(n521), .CO(n520), .S(product[61]) );
  FA_X1 U307 ( .A(n725), .B(n722), .CI(n522), .CO(n521), .S(product[60]) );
  FA_X1 U308 ( .A(n726), .B(n728), .CI(n523), .CO(n522), .S(product[59]) );
  FA_X1 U309 ( .A(n729), .B(n732), .CI(n524), .CO(n523), .S(product[58]) );
  FA_X1 U316 ( .A(n758), .B(n764), .CI(n529), .CO(n528), .S(product[53]) );
  FA_X1 U317 ( .A(n765), .B(n772), .CI(n530), .CO(n529), .S(product[52]) );
  FA_X1 U318 ( .A(n773), .B(n782), .CI(n531), .CO(n530), .S(product[51]) );
  FA_X1 U319 ( .A(n783), .B(n791), .CI(n532), .CO(n531), .S(product[50]) );
  FA_X1 U320 ( .A(n792), .B(n801), .CI(n533), .CO(n532), .S(product[49]) );
  FA_X1 U321 ( .A(n802), .B(n813), .CI(n534), .CO(n533), .S(product[48]) );
  FA_X1 U327 ( .A(n878), .B(n893), .CI(n540), .CO(n539), .S(product[42]) );
  FA_X1 U328 ( .A(n894), .B(n909), .CI(n541), .CO(n540), .S(product[41]) );
  FA_X1 U329 ( .A(n910), .B(n925), .CI(n542), .CO(n541), .S(product[40]) );
  FA_X1 U330 ( .A(n926), .B(n943), .CI(n543), .CO(n542), .S(product[39]) );
  FA_X1 U331 ( .A(n944), .B(n960), .CI(n544), .CO(n543), .S(product[38]) );
  FA_X1 U332 ( .A(n961), .B(n978), .CI(n545), .CO(n544), .S(product[37]) );
  FA_X1 U333 ( .A(n979), .B(n996), .CI(n546), .CO(n545), .S(product[36]) );
  FA_X1 U334 ( .A(n997), .B(n1014), .CI(n547), .CO(n546), .S(product[35]) );
  NAND2_X4 U337 ( .A1(n683), .A2(n549), .ZN(n486) );
  NOR2_X4 U339 ( .A1(n1015), .A2(n1032), .ZN(n548) );
  NAND2_X4 U340 ( .A1(n1015), .A2(n1032), .ZN(n549) );
  NAND2_X4 U345 ( .A1(n684), .A2(n554), .ZN(n487) );
  NOR2_X4 U347 ( .A1(n1033), .A2(n1050), .ZN(n553) );
  NAND2_X4 U348 ( .A1(n1033), .A2(n1050), .ZN(n554) );
  XOR2_X2 U349 ( .A(n558), .B(n488), .Z(product[32]) );
  NAND2_X4 U351 ( .A1(n685), .A2(n557), .ZN(n488) );
  NOR2_X4 U353 ( .A1(n1051), .A2(n1068), .ZN(n556) );
  NAND2_X4 U354 ( .A1(n1051), .A2(n1068), .ZN(n557) );
  AOI21_X4 U356 ( .B1(n563), .B2(n686), .A(n560), .ZN(n558) );
  NAND2_X4 U359 ( .A1(n686), .A2(n562), .ZN(n489) );
  NOR2_X4 U361 ( .A1(n1069), .A2(n1086), .ZN(n561) );
  NAND2_X4 U362 ( .A1(n1069), .A2(n1086), .ZN(n562) );
  NAND2_X4 U365 ( .A1(n687), .A2(n565), .ZN(n490) );
  NOR2_X4 U367 ( .A1(n1087), .A2(n1104), .ZN(n564) );
  NAND2_X4 U368 ( .A1(n1087), .A2(n1104), .ZN(n565) );
  NAND2_X4 U373 ( .A1(n688), .A2(n570), .ZN(n491) );
  NOR2_X4 U375 ( .A1(n1105), .A2(n1122), .ZN(n569) );
  NAND2_X4 U376 ( .A1(n1105), .A2(n1122), .ZN(n570) );
  XOR2_X2 U377 ( .A(n574), .B(n492), .Z(product[28]) );
  NAND2_X4 U379 ( .A1(n689), .A2(n573), .ZN(n492) );
  NOR2_X4 U381 ( .A1(n1123), .A2(n1140), .ZN(n572) );
  NAND2_X4 U382 ( .A1(n1123), .A2(n1140), .ZN(n573) );
  AOI21_X4 U384 ( .B1(n579), .B2(n690), .A(n576), .ZN(n574) );
  NAND2_X4 U387 ( .A1(n690), .A2(n578), .ZN(n493) );
  NOR2_X4 U389 ( .A1(n1141), .A2(n1158), .ZN(n577) );
  NAND2_X4 U390 ( .A1(n1141), .A2(n1158), .ZN(n578) );
  XOR2_X2 U391 ( .A(n582), .B(n494), .Z(product[26]) );
  NAND2_X4 U393 ( .A1(n691), .A2(n581), .ZN(n494) );
  NOR2_X4 U395 ( .A1(n1159), .A2(n1174), .ZN(n580) );
  NAND2_X4 U396 ( .A1(n1159), .A2(n1174), .ZN(n581) );
  AOI21_X4 U398 ( .B1(n587), .B2(n692), .A(n584), .ZN(n582) );
  NAND2_X4 U401 ( .A1(n692), .A2(n586), .ZN(n495) );
  NOR2_X4 U403 ( .A1(n1175), .A2(n1190), .ZN(n585) );
  NAND2_X4 U404 ( .A1(n1175), .A2(n1190), .ZN(n586) );
  NAND2_X4 U407 ( .A1(n693), .A2(n589), .ZN(n496) );
  NOR2_X4 U409 ( .A1(n1191), .A2(n1206), .ZN(n588) );
  NAND2_X4 U412 ( .A1(n1191), .A2(n1206), .ZN(n589) );
  AOI21_X4 U414 ( .B1(n595), .B2(n694), .A(n592), .ZN(n590) );
  NAND2_X4 U417 ( .A1(n694), .A2(n594), .ZN(n497) );
  NOR2_X4 U419 ( .A1(n1207), .A2(n1220), .ZN(n593) );
  NAND2_X4 U420 ( .A1(n1207), .A2(n1220), .ZN(n594) );
  NAND2_X4 U423 ( .A1(n695), .A2(n597), .ZN(n498) );
  NOR2_X4 U425 ( .A1(n1221), .A2(n1234), .ZN(n596) );
  NAND2_X4 U426 ( .A1(n1221), .A2(n1234), .ZN(n597) );
  AOI21_X4 U428 ( .B1(n603), .B2(n696), .A(n600), .ZN(n598) );
  NAND2_X4 U431 ( .A1(n696), .A2(n602), .ZN(n499) );
  NOR2_X4 U433 ( .A1(n1235), .A2(n1248), .ZN(n601) );
  NAND2_X4 U434 ( .A1(n1235), .A2(n1248), .ZN(n602) );
  XOR2_X2 U435 ( .A(n606), .B(n500), .Z(product[20]) );
  NAND2_X4 U437 ( .A1(n697), .A2(n605), .ZN(n500) );
  NOR2_X4 U439 ( .A1(n1249), .A2(n1260), .ZN(n604) );
  NAND2_X4 U440 ( .A1(n1249), .A2(n1260), .ZN(n605) );
  AOI21_X4 U442 ( .B1(n611), .B2(n698), .A(n608), .ZN(n606) );
  NAND2_X4 U445 ( .A1(n698), .A2(n610), .ZN(n501) );
  NOR2_X4 U447 ( .A1(n1261), .A2(n1272), .ZN(n609) );
  NAND2_X4 U448 ( .A1(n1261), .A2(n1272), .ZN(n610) );
  XOR2_X2 U449 ( .A(n614), .B(n502), .Z(product[18]) );
  NAND2_X4 U451 ( .A1(n699), .A2(n613), .ZN(n502) );
  NOR2_X4 U453 ( .A1(n1273), .A2(n1284), .ZN(n612) );
  NAND2_X4 U454 ( .A1(n1273), .A2(n1284), .ZN(n613) );
  AOI21_X4 U456 ( .B1(n619), .B2(n700), .A(n616), .ZN(n614) );
  NAND2_X4 U459 ( .A1(n700), .A2(n618), .ZN(n503) );
  NOR2_X4 U461 ( .A1(n1285), .A2(n1294), .ZN(n617) );
  NAND2_X4 U462 ( .A1(n1285), .A2(n1294), .ZN(n618) );
  XOR2_X2 U463 ( .A(n622), .B(n504), .Z(product[16]) );
  NAND2_X4 U465 ( .A1(n701), .A2(n621), .ZN(n504) );
  NOR2_X4 U467 ( .A1(n1295), .A2(n1304), .ZN(n620) );
  NAND2_X4 U468 ( .A1(n1295), .A2(n1304), .ZN(n621) );
  XNOR2_X2 U469 ( .A(n627), .B(n505), .ZN(product[15]) );
  AOI21_X4 U470 ( .B1(n627), .B2(n702), .A(n624), .ZN(n622) );
  NAND2_X4 U473 ( .A1(n702), .A2(n626), .ZN(n505) );
  NOR2_X4 U475 ( .A1(n1305), .A2(n1314), .ZN(n625) );
  NAND2_X4 U476 ( .A1(n1305), .A2(n1314), .ZN(n626) );
  XOR2_X2 U477 ( .A(n630), .B(n506), .Z(product[14]) );
  OAI21_X4 U478 ( .B1(n630), .B2(n628), .A(n629), .ZN(n627) );
  NAND2_X4 U479 ( .A1(n703), .A2(n629), .ZN(n506) );
  NOR2_X4 U481 ( .A1(n1315), .A2(n1322), .ZN(n628) );
  NAND2_X4 U482 ( .A1(n1315), .A2(n1322), .ZN(n629) );
  XNOR2_X2 U483 ( .A(n635), .B(n507), .ZN(product[13]) );
  AOI21_X4 U484 ( .B1(n635), .B2(n704), .A(n632), .ZN(n630) );
  NAND2_X4 U487 ( .A1(n704), .A2(n634), .ZN(n507) );
  NOR2_X4 U489 ( .A1(n1323), .A2(n1330), .ZN(n633) );
  NAND2_X4 U490 ( .A1(n1323), .A2(n1330), .ZN(n634) );
  XOR2_X2 U491 ( .A(n638), .B(n508), .Z(product[12]) );
  OAI21_X4 U492 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  NAND2_X4 U493 ( .A1(n705), .A2(n637), .ZN(n508) );
  NOR2_X4 U495 ( .A1(n1331), .A2(n1338), .ZN(n636) );
  NAND2_X4 U496 ( .A1(n1331), .A2(n1338), .ZN(n637) );
  AOI21_X4 U498 ( .B1(n643), .B2(n706), .A(n640), .ZN(n638) );
  NAND2_X4 U501 ( .A1(n706), .A2(n642), .ZN(n509) );
  NAND2_X4 U507 ( .A1(n707), .A2(n645), .ZN(n510) );
  NOR2_X4 U509 ( .A1(n1345), .A2(n1350), .ZN(n644) );
  NAND2_X4 U510 ( .A1(n1345), .A2(n1350), .ZN(n645) );
  AOI21_X4 U512 ( .B1(n651), .B2(n708), .A(n648), .ZN(n646) );
  NAND2_X4 U515 ( .A1(n708), .A2(n650), .ZN(n511) );
  XOR2_X2 U519 ( .A(n654), .B(n512), .Z(product[8]) );
  NAND2_X4 U521 ( .A1(n709), .A2(n653), .ZN(n512) );
  NOR2_X4 U523 ( .A1(n1357), .A2(n1360), .ZN(n652) );
  NAND2_X4 U524 ( .A1(n1357), .A2(n1360), .ZN(n653) );
  AOI21_X4 U526 ( .B1(n659), .B2(n710), .A(n656), .ZN(n654) );
  NAND2_X4 U529 ( .A1(n710), .A2(n658), .ZN(n513) );
  NOR2_X4 U531 ( .A1(n1361), .A2(n1364), .ZN(n657) );
  NAND2_X4 U532 ( .A1(n1361), .A2(n1364), .ZN(n658) );
  XOR2_X2 U533 ( .A(n514), .B(n662), .Z(product[6]) );
  NAND2_X4 U535 ( .A1(n711), .A2(n661), .ZN(n514) );
  NOR2_X4 U537 ( .A1(n1365), .A2(n2087), .ZN(n660) );
  NAND2_X4 U538 ( .A1(n1365), .A2(n2087), .ZN(n661) );
  XNOR2_X2 U539 ( .A(n515), .B(n667), .ZN(product[5]) );
  AOI21_X4 U540 ( .B1(n712), .B2(n667), .A(n664), .ZN(n662) );
  NAND2_X4 U543 ( .A1(n712), .A2(n666), .ZN(n515) );
  NOR2_X4 U545 ( .A1(n2088), .A2(n1369), .ZN(n665) );
  NAND2_X4 U546 ( .A1(n2088), .A2(n1369), .ZN(n666) );
  XOR2_X2 U547 ( .A(n516), .B(n670), .Z(product[4]) );
  OAI21_X4 U548 ( .B1(n670), .B2(n668), .A(n669), .ZN(n667) );
  NAND2_X4 U549 ( .A1(n713), .A2(n669), .ZN(n516) );
  NOR2_X4 U551 ( .A1(n1371), .A2(n2089), .ZN(n668) );
  NAND2_X4 U552 ( .A1(n1371), .A2(n2089), .ZN(n669) );
  XNOR2_X2 U553 ( .A(n517), .B(n675), .ZN(product[3]) );
  AOI21_X4 U554 ( .B1(n675), .B2(n714), .A(n672), .ZN(n670) );
  NAND2_X4 U557 ( .A1(n714), .A2(n674), .ZN(n517) );
  XOR2_X2 U561 ( .A(n676), .B(n677), .Z(product[2]) );
  NOR2_X4 U562 ( .A1(n676), .A2(n677), .ZN(n675) );
  XNOR2_X2 U564 ( .A(n679), .B(n680), .ZN(product[1]) );
  NAND2_X4 U565 ( .A1(n678), .A2(n680), .ZN(n677) );
  NAND2_X4 U570 ( .A1(n715), .A2(n682), .ZN(n518) );
  NOR2_X4 U572 ( .A1(n2093), .A2(n262), .ZN(n681) );
  NAND2_X4 U573 ( .A1(n2093), .A2(n262), .ZN(n682) );
  FA_X1 U576 ( .A(n1721), .B(n1745), .CI(n723), .CO(n719), .S(n720) );
  FA_X1 U577 ( .A(n727), .B(n1722), .CI(n1746), .CO(n721), .S(n722) );
  FA_X1 U579 ( .A(n1747), .B(n727), .CI(n730), .CO(n725), .S(n726) );
  FA_X1 U581 ( .A(n734), .B(n1748), .CI(n731), .CO(n728), .S(n729) );
  FA_X1 U582 ( .A(n736), .B(n1779), .CI(n1723), .CO(n730), .S(n731) );
  FA_X1 U583 ( .A(n740), .B(n1749), .CI(n735), .CO(n732), .S(n733) );
  FA_X1 U584 ( .A(n742), .B(n1724), .CI(n1780), .CO(n734), .S(n735) );
  FA_X1 U586 ( .A(n741), .B(n747), .CI(n745), .CO(n738), .S(n739) );
  FA_X1 U587 ( .A(n1781), .B(n742), .CI(n1750), .CO(n740), .S(n741) );
  FA_X1 U589 ( .A(n751), .B(n748), .CI(n746), .CO(n743), .S(n744) );
  FA_X1 U590 ( .A(n1751), .B(n1782), .CI(n753), .CO(n745), .S(n746) );
  FA_X1 U591 ( .A(n755), .B(n1814), .CI(n1725), .CO(n747), .S(n748) );
  FA_X1 U592 ( .A(n759), .B(n754), .CI(n752), .CO(n749), .S(n750) );
  FA_X1 U593 ( .A(n1752), .B(n1783), .CI(n761), .CO(n751), .S(n752) );
  FA_X1 U594 ( .A(n763), .B(n1726), .CI(n1815), .CO(n753), .S(n754) );
  FA_X1 U596 ( .A(n766), .B(n762), .CI(n760), .CO(n757), .S(n758) );
  FA_X1 U597 ( .A(n770), .B(n1753), .CI(n768), .CO(n759), .S(n760) );
  FA_X1 U598 ( .A(n1816), .B(n763), .CI(n1784), .CO(n761), .S(n762) );
  FA_X1 U600 ( .A(n774), .B(n769), .CI(n767), .CO(n764), .S(n765) );
  FA_X1 U601 ( .A(n771), .B(n778), .CI(n776), .CO(n766), .S(n767) );
  FA_X1 U602 ( .A(n1785), .B(n1754), .CI(n1817), .CO(n768), .S(n769) );
  FA_X1 U603 ( .A(n780), .B(n1849), .CI(n1727), .CO(n770), .S(n771) );
  FA_X1 U604 ( .A(n784), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U605 ( .A(n779), .B(n788), .CI(n786), .CO(n774), .S(n775) );
  FA_X1 U606 ( .A(n1786), .B(n1755), .CI(n1818), .CO(n776), .S(n777) );
  FA_X1 U607 ( .A(n790), .B(n1728), .CI(n1850), .CO(n778), .S(n779) );
  FA_X1 U609 ( .A(n793), .B(n787), .CI(n785), .CO(n782), .S(n783) );
  FA_X1 U610 ( .A(n789), .B(n797), .CI(n795), .CO(n784), .S(n785) );
  FA_X1 U611 ( .A(n1787), .B(n1819), .CI(n799), .CO(n786), .S(n787) );
  FA_X1 U612 ( .A(n1851), .B(n790), .CI(n1756), .CO(n788), .S(n789) );
  FA_X1 U614 ( .A(n803), .B(n796), .CI(n794), .CO(n791), .S(n792) );
  FA_X1 U615 ( .A(n798), .B(n807), .CI(n805), .CO(n793), .S(n794) );
  FA_X1 U616 ( .A(n809), .B(n1820), .CI(n800), .CO(n795), .S(n796) );
  FA_X1 U617 ( .A(n1852), .B(n1757), .CI(n1788), .CO(n797), .S(n798) );
  FA_X1 U618 ( .A(n811), .B(n1884), .CI(n1729), .CO(n799), .S(n800) );
  FA_X1 U619 ( .A(n815), .B(n806), .CI(n804), .CO(n801), .S(n802) );
  FA_X1 U620 ( .A(n808), .B(n819), .CI(n817), .CO(n803), .S(n804) );
  FA_X1 U621 ( .A(n821), .B(n1758), .CI(n810), .CO(n805), .S(n806) );
  FA_X1 U622 ( .A(n1853), .B(n1789), .CI(n1821), .CO(n807), .S(n808) );
  FA_X1 U623 ( .A(n823), .B(n1730), .CI(n1885), .CO(n809), .S(n810) );
  FA_X1 U625 ( .A(n826), .B(n818), .CI(n816), .CO(n813), .S(n814) );
  FA_X1 U626 ( .A(n820), .B(n822), .CI(n828), .CO(n815), .S(n816) );
  FA_X1 U627 ( .A(n832), .B(n1759), .CI(n830), .CO(n817), .S(n818) );
  FA_X1 U628 ( .A(n1822), .B(n1790), .CI(n1854), .CO(n819), .S(n820) );
  FA_X1 U629 ( .A(n834), .B(n823), .CI(n1886), .CO(n821), .S(n822) );
  FA_X1 U631 ( .A(n838), .B(n829), .CI(n827), .CO(n824), .S(n825) );
  FA_X1 U632 ( .A(n842), .B(n833), .CI(n840), .CO(n826), .S(n827) );
  FA_X1 U633 ( .A(n844), .B(n846), .CI(n831), .CO(n828), .S(n829) );
  FA_X1 U634 ( .A(n1823), .B(n1760), .CI(n1887), .CO(n830), .S(n831) );
  FA_X1 U635 ( .A(n1855), .B(n1791), .CI(n835), .CO(n832), .S(n833) );
  FA_X1 U636 ( .A(n848), .B(n1919), .CI(n1731), .CO(n834), .S(n835) );
  FA_X1 U637 ( .A(n852), .B(n841), .CI(n839), .CO(n836), .S(n837) );
  FA_X1 U638 ( .A(n843), .B(n856), .CI(n854), .CO(n838), .S(n839) );
  FA_X1 U639 ( .A(n858), .B(n847), .CI(n845), .CO(n840), .S(n841) );
  FA_X1 U640 ( .A(n1761), .B(n1824), .CI(n860), .CO(n842), .S(n843) );
  FA_X1 U641 ( .A(n1888), .B(n1792), .CI(n1856), .CO(n844), .S(n845) );
  FA_X1 U642 ( .A(n1732), .B(n862), .CI(n1920), .CO(n846), .S(n847) );
  FA_X1 U644 ( .A(n865), .B(n855), .CI(n853), .CO(n850), .S(n851) );
  FA_X1 U645 ( .A(n857), .B(n869), .CI(n867), .CO(n852), .S(n853) );
  FA_X1 U646 ( .A(n861), .B(n871), .CI(n859), .CO(n854), .S(n855) );
  FA_X1 U647 ( .A(n1857), .B(n1762), .CI(n873), .CO(n856), .S(n857) );
  FA_X1 U648 ( .A(n1889), .B(n1793), .CI(n875), .CO(n858), .S(n859) );
  FA_X1 U649 ( .A(n1921), .B(n862), .CI(n1825), .CO(n860), .S(n861) );
  FA_X1 U651 ( .A(n879), .B(n868), .CI(n866), .CO(n863), .S(n864) );
  FA_X1 U652 ( .A(n870), .B(n883), .CI(n881), .CO(n865), .S(n866) );
  FA_X1 U653 ( .A(n874), .B(n885), .CI(n872), .CO(n867), .S(n868) );
  FA_X1 U654 ( .A(n889), .B(n876), .CI(n887), .CO(n869), .S(n870) );
  FA_X1 U655 ( .A(n1858), .B(n1922), .CI(n1890), .CO(n871), .S(n872) );
  FA_X1 U656 ( .A(n1826), .B(n1763), .CI(n1794), .CO(n873), .S(n874) );
  FA_X1 U657 ( .A(n891), .B(n3224), .CI(n1733), .CO(n875), .S(n876) );
  FA_X1 U658 ( .A(n895), .B(n882), .CI(n880), .CO(n877), .S(n878) );
  FA_X1 U659 ( .A(n884), .B(n899), .CI(n897), .CO(n879), .S(n880) );
  FA_X1 U660 ( .A(n888), .B(n901), .CI(n886), .CO(n881), .S(n882) );
  FA_X1 U661 ( .A(n890), .B(n905), .CI(n903), .CO(n883), .S(n884) );
  FA_X1 U662 ( .A(n1891), .B(n1859), .CI(n1923), .CO(n885), .S(n886) );
  FA_X1 U663 ( .A(n1827), .B(n1764), .CI(n1795), .CO(n887), .S(n888) );
  FA_X1 U664 ( .A(n907), .B(n892), .CI(n1955), .CO(n889), .S(n890) );
  FA_X1 U666 ( .A(n911), .B(n898), .CI(n896), .CO(n893), .S(n894) );
  FA_X1 U667 ( .A(n900), .B(n915), .CI(n913), .CO(n895), .S(n896) );
  FA_X1 U668 ( .A(n904), .B(n917), .CI(n902), .CO(n897), .S(n898) );
  FA_X1 U669 ( .A(n921), .B(n906), .CI(n919), .CO(n899), .S(n900) );
  FA_X1 U670 ( .A(n1892), .B(n1796), .CI(n1924), .CO(n901), .S(n902) );
  FA_X1 U671 ( .A(n1828), .B(n1956), .CI(n1860), .CO(n903), .S(n904) );
  FA_X1 U672 ( .A(n908), .B(n1734), .CI(n923), .CO(n905), .S(n906) );
  FA_X1 U674 ( .A(n927), .B(n914), .CI(n912), .CO(n909), .S(n910) );
  FA_X1 U675 ( .A(n916), .B(n931), .CI(n929), .CO(n911), .S(n912) );
  FA_X1 U676 ( .A(n920), .B(n933), .CI(n918), .CO(n913), .S(n914) );
  FA_X1 U677 ( .A(n935), .B(n937), .CI(n922), .CO(n915), .S(n916) );
  FA_X1 U678 ( .A(n1893), .B(n1829), .CI(n1957), .CO(n917), .S(n918) );
  FA_X1 U679 ( .A(n1925), .B(n1861), .CI(n939), .CO(n919), .S(n920) );
  FA_X1 U680 ( .A(n1765), .B(n1797), .CI(n924), .CO(n921), .S(n922) );
  FA_X1 U681 ( .A(n941), .B(n3229), .CI(n1735), .CO(n923), .S(n924) );
  FA_X1 U682 ( .A(n945), .B(n930), .CI(n928), .CO(n925), .S(n926) );
  FA_X1 U683 ( .A(n932), .B(n949), .CI(n947), .CO(n927), .S(n928) );
  FA_X1 U684 ( .A(n951), .B(n936), .CI(n934), .CO(n929), .S(n930) );
  FA_X1 U685 ( .A(n953), .B(n955), .CI(n938), .CO(n931), .S(n932) );
  FA_X1 U686 ( .A(n957), .B(n1894), .CI(n940), .CO(n933), .S(n934) );
  FA_X1 U687 ( .A(n1926), .B(n1830), .CI(n1958), .CO(n935), .S(n936) );
  FA_X1 U688 ( .A(n1798), .B(n1990), .CI(n1862), .CO(n937), .S(n938) );
  FA_X1 U689 ( .A(n1736), .B(n959), .CI(n1766), .CO(n939), .S(n940) );
  FA_X1 U691 ( .A(n962), .B(n948), .CI(n946), .CO(n943), .S(n944) );
  FA_X1 U692 ( .A(n950), .B(n966), .CI(n964), .CO(n945), .S(n946) );
  FA_X1 U693 ( .A(n968), .B(n954), .CI(n952), .CO(n947), .S(n948) );
  FA_X1 U694 ( .A(n970), .B(n972), .CI(n956), .CO(n949), .S(n950) );
  FA_X1 U695 ( .A(n974), .B(n1895), .CI(n958), .CO(n951), .S(n952) );
  FA_X1 U696 ( .A(n1927), .B(n1831), .CI(n1959), .CO(n953), .S(n954) );
  FA_X1 U697 ( .A(n1767), .B(n1991), .CI(n1863), .CO(n955), .S(n956) );
  FA_X1 U698 ( .A(n1799), .B(n959), .CI(n976), .CO(n957), .S(n958) );
  FA_X1 U700 ( .A(n980), .B(n965), .CI(n963), .CO(n960), .S(n961) );
  FA_X1 U701 ( .A(n967), .B(n969), .CI(n982), .CO(n962), .S(n963) );
  FA_X1 U702 ( .A(n986), .B(n971), .CI(n984), .CO(n964), .S(n965) );
  FA_X1 U703 ( .A(n975), .B(n988), .CI(n973), .CO(n966), .S(n967) );
  FA_X1 U704 ( .A(n992), .B(n1960), .CI(n990), .CO(n968), .S(n969) );
  FA_X1 U705 ( .A(n1928), .B(n1992), .CI(n994), .CO(n970), .S(n971) );
  FA_X1 U706 ( .A(n1896), .B(n977), .CI(n1864), .CO(n972), .S(n973) );
  FA_X1 U707 ( .A(n1832), .B(n1768), .CI(n1800), .CO(n974), .S(n975) );
  FA_X1 U708 ( .A(n3232), .B(n2059), .CI(n1737), .CO(n976), .S(n977) );
  FA_X1 U709 ( .A(n998), .B(n983), .CI(n981), .CO(n978), .S(n979) );
  FA_X1 U710 ( .A(n985), .B(n987), .CI(n1000), .CO(n980), .S(n981) );
  FA_X1 U711 ( .A(n1004), .B(n989), .CI(n1002), .CO(n982), .S(n983) );
  FA_X1 U712 ( .A(n993), .B(n1006), .CI(n991), .CO(n984), .S(n985) );
  FA_X1 U713 ( .A(n1010), .B(n995), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U714 ( .A(n1865), .B(n1929), .CI(n1961), .CO(n988), .S(n989) );
  FA_X1 U715 ( .A(n1897), .B(n1012), .CI(n1993), .CO(n990), .S(n991) );
  FA_X1 U716 ( .A(n2025), .B(n1769), .CI(n1833), .CO(n992), .S(n993) );
  FA_X1 U717 ( .A(n1738), .B(n262), .CI(n1801), .CO(n994), .S(n995) );
  FA_X1 U718 ( .A(n1016), .B(n1001), .CI(n999), .CO(n996), .S(n997) );
  FA_X1 U719 ( .A(n1003), .B(n1005), .CI(n1018), .CO(n998), .S(n999) );
  FA_X1 U720 ( .A(n1022), .B(n1009), .CI(n1020), .CO(n1000), .S(n1001) );
  FA_X1 U721 ( .A(n1011), .B(n1024), .CI(n1007), .CO(n1002), .S(n1003) );
  FA_X1 U722 ( .A(n1028), .B(n1013), .CI(n1026), .CO(n1004), .S(n1005) );
  FA_X1 U723 ( .A(n1866), .B(n1930), .CI(n1962), .CO(n1006), .S(n1007) );
  FA_X1 U724 ( .A(n1994), .B(n1898), .CI(n1030), .CO(n1008), .S(n1009) );
  FA_X1 U725 ( .A(n2026), .B(n1834), .CI(n1802), .CO(n1010), .S(n1011) );
  FA_X1 U726 ( .A(n1739), .B(n262), .CI(n1770), .CO(n1012), .S(n1013) );
  FA_X1 U727 ( .A(n1034), .B(n1019), .CI(n1017), .CO(n1014), .S(n1015) );
  FA_X1 U728 ( .A(n1021), .B(n1023), .CI(n1036), .CO(n1016), .S(n1017) );
  FA_X1 U729 ( .A(n1040), .B(n1027), .CI(n1038), .CO(n1018), .S(n1019) );
  FA_X1 U730 ( .A(n1029), .B(n1042), .CI(n1025), .CO(n1020), .S(n1021) );
  FA_X1 U731 ( .A(n1046), .B(n1031), .CI(n1044), .CO(n1022), .S(n1023) );
  FA_X1 U732 ( .A(n1963), .B(n1899), .CI(n1995), .CO(n1024), .S(n1025) );
  FA_X1 U733 ( .A(n2027), .B(n1931), .CI(n1048), .CO(n1026), .S(n1027) );
  FA_X1 U734 ( .A(n1867), .B(n1803), .CI(n1835), .CO(n1028), .S(n1029) );
  FA_X1 U735 ( .A(n1740), .B(n262), .CI(n1771), .CO(n1030), .S(n1031) );
  FA_X1 U736 ( .A(n1052), .B(n1037), .CI(n1035), .CO(n1032), .S(n1033) );
  FA_X1 U737 ( .A(n1039), .B(n1041), .CI(n1054), .CO(n1034), .S(n1035) );
  FA_X1 U738 ( .A(n1058), .B(n1045), .CI(n1056), .CO(n1036), .S(n1037) );
  FA_X1 U739 ( .A(n1047), .B(n1060), .CI(n1043), .CO(n1038), .S(n1039) );
  FA_X1 U740 ( .A(n1064), .B(n1049), .CI(n1062), .CO(n1040), .S(n1041) );
  FA_X1 U741 ( .A(n1900), .B(n1964), .CI(n1066), .CO(n1042), .S(n1043) );
  FA_X1 U742 ( .A(n2028), .B(n1932), .CI(n1996), .CO(n1044), .S(n1045) );
  FA_X1 U743 ( .A(n2060), .B(n1836), .CI(n1868), .CO(n1046), .S(n1047) );
  FA_X1 U744 ( .A(n1772), .B(n1741), .CI(n1804), .CO(n1048), .S(n1049) );
  FA_X1 U745 ( .A(n1070), .B(n1055), .CI(n1053), .CO(n1050), .S(n1051) );
  FA_X1 U746 ( .A(n1057), .B(n1059), .CI(n1072), .CO(n1052), .S(n1053) );
  FA_X1 U747 ( .A(n1076), .B(n1063), .CI(n1074), .CO(n1054), .S(n1055) );
  FA_X1 U748 ( .A(n1065), .B(n1078), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U749 ( .A(n1067), .B(n1082), .CI(n1080), .CO(n1058), .S(n1059) );
  FA_X1 U750 ( .A(n1933), .B(n1965), .CI(n1997), .CO(n1060), .S(n1061) );
  FA_X1 U751 ( .A(n2029), .B(n1901), .CI(n1084), .CO(n1062), .S(n1063) );
  FA_X1 U752 ( .A(n2061), .B(n1869), .CI(n1837), .CO(n1064), .S(n1065) );
  FA_X1 U753 ( .A(n1773), .B(n1742), .CI(n1805), .CO(n1066), .S(n1067) );
  FA_X1 U754 ( .A(n1088), .B(n1073), .CI(n1071), .CO(n1068), .S(n1069) );
  FA_X1 U755 ( .A(n1075), .B(n1092), .CI(n1090), .CO(n1070), .S(n1071) );
  FA_X1 U756 ( .A(n1079), .B(n1094), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U757 ( .A(n1096), .B(n1098), .CI(n1081), .CO(n1074), .S(n1075) );
  FA_X1 U758 ( .A(n1085), .B(n1100), .CI(n1083), .CO(n1076), .S(n1077) );
  FA_X1 U759 ( .A(n1998), .B(n2062), .CI(n2030), .CO(n1078), .S(n1079) );
  FA_X1 U760 ( .A(n1966), .B(n1870), .CI(n1934), .CO(n1080), .S(n1081) );
  FA_X1 U761 ( .A(n1102), .B(n1838), .CI(n1902), .CO(n1082), .S(n1083) );
  FA_X1 U762 ( .A(n1774), .B(n1743), .CI(n1806), .CO(n1084), .S(n1085) );
  FA_X1 U763 ( .A(n1106), .B(n1091), .CI(n1089), .CO(n1086), .S(n1087) );
  FA_X1 U764 ( .A(n1108), .B(n1110), .CI(n1093), .CO(n1088), .S(n1089) );
  FA_X1 U765 ( .A(n1097), .B(n1099), .CI(n1095), .CO(n1090), .S(n1091) );
  FA_X1 U766 ( .A(n1114), .B(n1116), .CI(n1112), .CO(n1092), .S(n1093) );
  FA_X1 U767 ( .A(n1118), .B(n1999), .CI(n1101), .CO(n1094), .S(n1095) );
  FA_X1 U768 ( .A(n2063), .B(n1935), .CI(n2031), .CO(n1096), .S(n1097) );
  FA_X1 U769 ( .A(n1903), .B(n1103), .CI(n1967), .CO(n1098), .S(n1099) );
  FA_X1 U770 ( .A(n1871), .B(n1807), .CI(n1839), .CO(n1100), .S(n1101) );
  FA_X1 U771 ( .A(n1775), .B(n1744), .CI(n1120), .CO(n1102), .S(n1103) );
  FA_X1 U772 ( .A(n1124), .B(n1109), .CI(n1107), .CO(n1104), .S(n1105) );
  FA_X1 U773 ( .A(n1126), .B(n1128), .CI(n1111), .CO(n1106), .S(n1107) );
  FA_X1 U774 ( .A(n1115), .B(n1117), .CI(n1113), .CO(n1108), .S(n1109) );
  FA_X1 U775 ( .A(n1132), .B(n1119), .CI(n1130), .CO(n1110), .S(n1111) );
  FA_X1 U776 ( .A(n2064), .B(n2000), .CI(n1134), .CO(n1112), .S(n1113) );
  FA_X1 U777 ( .A(n2032), .B(n1936), .CI(n1136), .CO(n1114), .S(n1115) );
  FA_X1 U778 ( .A(n1872), .B(n1904), .CI(n1968), .CO(n1116), .S(n1117) );
  FA_X1 U779 ( .A(n1808), .B(n1121), .CI(n1840), .CO(n1118), .S(n1119) );
  HA_X1 U780 ( .A(n1776), .B(n1138), .CO(n1120), .S(n1121) );
  FA_X1 U781 ( .A(n1142), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U782 ( .A(n1129), .B(n1146), .CI(n1144), .CO(n1124), .S(n1125) );
  FA_X1 U783 ( .A(n1133), .B(n1148), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U784 ( .A(n1135), .B(n1137), .CI(n1150), .CO(n1128), .S(n1129) );
  FA_X1 U785 ( .A(n2033), .B(n2065), .CI(n1152), .CO(n1130), .S(n1131) );
  FA_X1 U786 ( .A(n2001), .B(n1905), .CI(n1969), .CO(n1132), .S(n1133) );
  FA_X1 U787 ( .A(n1154), .B(n1873), .CI(n1937), .CO(n1134), .S(n1135) );
  FA_X1 U788 ( .A(n1139), .B(n1809), .CI(n1841), .CO(n1136), .S(n1137) );
  HA_X1 U789 ( .A(n1156), .B(n1777), .CO(n1138), .S(n1139) );
  FA_X1 U790 ( .A(n1160), .B(n1145), .CI(n1143), .CO(n1140), .S(n1141) );
  FA_X1 U791 ( .A(n1147), .B(n1149), .CI(n1162), .CO(n1142), .S(n1143) );
  FA_X1 U792 ( .A(n1164), .B(n1166), .CI(n1151), .CO(n1144), .S(n1145) );
  FA_X1 U793 ( .A(n1153), .B(n2002), .CI(n1168), .CO(n1146), .S(n1147) );
  FA_X1 U794 ( .A(n1170), .B(n2034), .CI(n2066), .CO(n1148), .S(n1149) );
  FA_X1 U795 ( .A(n1938), .B(n1155), .CI(n1970), .CO(n1150), .S(n1151) );
  FA_X1 U796 ( .A(n1874), .B(n1842), .CI(n1906), .CO(n1152), .S(n1153) );
  FA_X1 U797 ( .A(n1810), .B(n1157), .CI(n1172), .CO(n1154), .S(n1155) );
  HA_X1 U798 ( .A(n289), .B(n1778), .CO(n1156), .S(n1157) );
  FA_X1 U799 ( .A(n1176), .B(n1163), .CI(n1161), .CO(n1158), .S(n1159) );
  FA_X1 U800 ( .A(n1165), .B(n1167), .CI(n1178), .CO(n1160), .S(n1161) );
  FA_X1 U801 ( .A(n1169), .B(n1182), .CI(n1180), .CO(n1162), .S(n1163) );
  FA_X1 U802 ( .A(n1184), .B(n2003), .CI(n1171), .CO(n1164), .S(n1165) );
  FA_X1 U803 ( .A(n2067), .B(n2035), .CI(n1186), .CO(n1166), .S(n1167) );
  FA_X1 U804 ( .A(n1907), .B(n1939), .CI(n1971), .CO(n1168), .S(n1169) );
  FA_X1 U805 ( .A(n1843), .B(n1173), .CI(n1875), .CO(n1170), .S(n1171) );
  HA_X1 U806 ( .A(n1811), .B(n1188), .CO(n1172), .S(n1173) );
  FA_X1 U807 ( .A(n1192), .B(n1179), .CI(n1177), .CO(n1174), .S(n1175) );
  FA_X1 U808 ( .A(n1181), .B(n1183), .CI(n1194), .CO(n1176), .S(n1177) );
  FA_X1 U809 ( .A(n1198), .B(n1185), .CI(n1196), .CO(n1178), .S(n1179) );
  FA_X1 U810 ( .A(n1200), .B(n2068), .CI(n1187), .CO(n1180), .S(n1181) );
  FA_X1 U811 ( .A(n2004), .B(n1940), .CI(n2036), .CO(n1182), .S(n1183) );
  FA_X1 U812 ( .A(n1202), .B(n1908), .CI(n1972), .CO(n1184), .S(n1185) );
  FA_X1 U813 ( .A(n1189), .B(n1844), .CI(n1876), .CO(n1186), .S(n1187) );
  HA_X1 U814 ( .A(n1204), .B(n1812), .CO(n1188), .S(n1189) );
  FA_X1 U815 ( .A(n1208), .B(n1195), .CI(n1193), .CO(n1190), .S(n1191) );
  FA_X1 U816 ( .A(n1197), .B(n1199), .CI(n1210), .CO(n1192), .S(n1193) );
  FA_X1 U817 ( .A(n1214), .B(n1201), .CI(n1212), .CO(n1194), .S(n1195) );
  FA_X1 U818 ( .A(n2037), .B(n2069), .CI(n1216), .CO(n1196), .S(n1197) );
  FA_X1 U819 ( .A(n1973), .B(n1203), .CI(n2005), .CO(n1198), .S(n1199) );
  FA_X1 U820 ( .A(n1941), .B(n1877), .CI(n1909), .CO(n1200), .S(n1201) );
  FA_X1 U821 ( .A(n1845), .B(n1205), .CI(n1218), .CO(n1202), .S(n1203) );
  HA_X1 U822 ( .A(n286), .B(n1813), .CO(n1204), .S(n1205) );
  FA_X1 U823 ( .A(n1222), .B(n1211), .CI(n1209), .CO(n1206), .S(n1207) );
  FA_X1 U824 ( .A(n1213), .B(n1215), .CI(n1224), .CO(n1208), .S(n1209) );
  FA_X1 U825 ( .A(n1217), .B(n1228), .CI(n1226), .CO(n1210), .S(n1211) );
  FA_X1 U826 ( .A(n2038), .B(n2070), .CI(n1230), .CO(n1212), .S(n1213) );
  FA_X1 U827 ( .A(n1942), .B(n1974), .CI(n2006), .CO(n1214), .S(n1215) );
  FA_X1 U828 ( .A(n1878), .B(n1219), .CI(n1910), .CO(n1216), .S(n1217) );
  HA_X1 U829 ( .A(n1846), .B(n1232), .CO(n1218), .S(n1219) );
  FA_X1 U830 ( .A(n1236), .B(n1225), .CI(n1223), .CO(n1220), .S(n1221) );
  FA_X1 U831 ( .A(n1227), .B(n1240), .CI(n1238), .CO(n1222), .S(n1223) );
  FA_X1 U832 ( .A(n1231), .B(n1242), .CI(n1229), .CO(n1224), .S(n1225) );
  FA_X1 U833 ( .A(n2071), .B(n1975), .CI(n2039), .CO(n1226), .S(n1227) );
  FA_X1 U834 ( .A(n1244), .B(n1943), .CI(n2007), .CO(n1228), .S(n1229) );
  FA_X1 U835 ( .A(n1233), .B(n1879), .CI(n1911), .CO(n1230), .S(n1231) );
  HA_X1 U836 ( .A(n1246), .B(n1847), .CO(n1232), .S(n1233) );
  FA_X1 U837 ( .A(n1250), .B(n1239), .CI(n1237), .CO(n1234), .S(n1235) );
  FA_X1 U838 ( .A(n1252), .B(n1254), .CI(n1241), .CO(n1236), .S(n1237) );
  FA_X1 U839 ( .A(n1256), .B(n2040), .CI(n1243), .CO(n1238), .S(n1239) );
  FA_X1 U840 ( .A(n2008), .B(n1245), .CI(n2072), .CO(n1240), .S(n1241) );
  FA_X1 U841 ( .A(n1944), .B(n1912), .CI(n1976), .CO(n1242), .S(n1243) );
  FA_X1 U842 ( .A(n1880), .B(n1247), .CI(n1258), .CO(n1244), .S(n1245) );
  HA_X1 U843 ( .A(n283), .B(n1848), .CO(n1246), .S(n1247) );
  FA_X1 U844 ( .A(n1262), .B(n1253), .CI(n1251), .CO(n1248), .S(n1249) );
  FA_X1 U845 ( .A(n1264), .B(n1257), .CI(n1255), .CO(n1250), .S(n1251) );
  FA_X1 U846 ( .A(n1268), .B(n2041), .CI(n1266), .CO(n1252), .S(n1253) );
  FA_X1 U847 ( .A(n1977), .B(n2009), .CI(n2073), .CO(n1254), .S(n1255) );
  FA_X1 U848 ( .A(n1913), .B(n1259), .CI(n1945), .CO(n1256), .S(n1257) );
  HA_X1 U849 ( .A(n1881), .B(n1270), .CO(n1258), .S(n1259) );
  FA_X1 U850 ( .A(n1274), .B(n1265), .CI(n1263), .CO(n1260), .S(n1261) );
  FA_X1 U851 ( .A(n1267), .B(n1269), .CI(n1276), .CO(n1262), .S(n1263) );
  FA_X1 U852 ( .A(n2074), .B(n2010), .CI(n1278), .CO(n1264), .S(n1265) );
  FA_X1 U853 ( .A(n1280), .B(n1978), .CI(n2042), .CO(n1266), .S(n1267) );
  FA_X1 U854 ( .A(n1271), .B(n1914), .CI(n1946), .CO(n1268), .S(n1269) );
  HA_X1 U855 ( .A(n1282), .B(n1882), .CO(n1270), .S(n1271) );
  FA_X1 U856 ( .A(n1277), .B(n1286), .CI(n1275), .CO(n1272), .S(n1273) );
  FA_X1 U857 ( .A(n1279), .B(n1290), .CI(n1288), .CO(n1274), .S(n1275) );
  FA_X1 U858 ( .A(n2043), .B(n1281), .CI(n2075), .CO(n1276), .S(n1277) );
  FA_X1 U859 ( .A(n2011), .B(n1947), .CI(n1979), .CO(n1278), .S(n1279) );
  FA_X1 U860 ( .A(n1915), .B(n1283), .CI(n1292), .CO(n1280), .S(n1281) );
  HA_X1 U861 ( .A(n280), .B(n1883), .CO(n1282), .S(n1283) );
  FA_X1 U862 ( .A(n1296), .B(n1289), .CI(n1287), .CO(n1284), .S(n1285) );
  FA_X1 U863 ( .A(n1298), .B(n1300), .CI(n1291), .CO(n1286), .S(n1287) );
  FA_X1 U864 ( .A(n2012), .B(n2044), .CI(n2076), .CO(n1288), .S(n1289) );
  FA_X1 U865 ( .A(n1948), .B(n1293), .CI(n1980), .CO(n1290), .S(n1291) );
  HA_X1 U866 ( .A(n1916), .B(n1302), .CO(n1292), .S(n1293) );
  FA_X1 U867 ( .A(n1306), .B(n1299), .CI(n1297), .CO(n1294), .S(n1295) );
  FA_X1 U868 ( .A(n1308), .B(n2045), .CI(n1301), .CO(n1296), .S(n1297) );
  FA_X1 U869 ( .A(n1310), .B(n2013), .CI(n2077), .CO(n1298), .S(n1299) );
  FA_X1 U870 ( .A(n1303), .B(n1949), .CI(n1981), .CO(n1300), .S(n1301) );
  HA_X1 U871 ( .A(n1312), .B(n1917), .CO(n1302), .S(n1303) );
  FA_X1 U872 ( .A(n1316), .B(n1309), .CI(n1307), .CO(n1304), .S(n1305) );
  FA_X1 U873 ( .A(n2078), .B(n1311), .CI(n1318), .CO(n1306), .S(n1307) );
  FA_X1 U874 ( .A(n2046), .B(n1982), .CI(n2014), .CO(n1308), .S(n1309) );
  FA_X1 U875 ( .A(n1950), .B(n1313), .CI(n1320), .CO(n1310), .S(n1311) );
  HA_X1 U876 ( .A(n277), .B(n1918), .CO(n1312), .S(n1313) );
  FA_X1 U877 ( .A(n1324), .B(n1319), .CI(n1317), .CO(n1314), .S(n1315) );
  FA_X1 U878 ( .A(n2047), .B(n2079), .CI(n1326), .CO(n1316), .S(n1317) );
  FA_X1 U879 ( .A(n1983), .B(n1321), .CI(n2015), .CO(n1318), .S(n1319) );
  HA_X1 U880 ( .A(n1951), .B(n1328), .CO(n1320), .S(n1321) );
  FA_X1 U881 ( .A(n1327), .B(n1332), .CI(n1325), .CO(n1322), .S(n1323) );
  FA_X1 U882 ( .A(n1334), .B(n2048), .CI(n2080), .CO(n1324), .S(n1325) );
  FA_X1 U883 ( .A(n1329), .B(n1984), .CI(n2016), .CO(n1326), .S(n1327) );
  HA_X1 U884 ( .A(n1336), .B(n1952), .CO(n1328), .S(n1329) );
  FA_X1 U885 ( .A(n1340), .B(n1335), .CI(n1333), .CO(n1330), .S(n1331) );
  FA_X1 U886 ( .A(n2081), .B(n2017), .CI(n2049), .CO(n1332), .S(n1333) );
  FA_X1 U887 ( .A(n1985), .B(n1337), .CI(n1342), .CO(n1334), .S(n1335) );
  HA_X1 U888 ( .A(n274), .B(n1953), .CO(n1336), .S(n1337) );
  FA_X1 U889 ( .A(n1346), .B(n2082), .CI(n1341), .CO(n1338), .S(n1339) );
  FA_X1 U890 ( .A(n2018), .B(n1343), .CI(n2050), .CO(n1340), .S(n1341) );
  HA_X1 U891 ( .A(n1986), .B(n1348), .CO(n1342), .S(n1343) );
  FA_X1 U892 ( .A(n1352), .B(n2083), .CI(n1347), .CO(n1344), .S(n1345) );
  FA_X1 U893 ( .A(n1349), .B(n2019), .CI(n2051), .CO(n1346), .S(n1347) );
  HA_X1 U894 ( .A(n1354), .B(n1987), .CO(n1348), .S(n1349) );
  FA_X1 U895 ( .A(n2084), .B(n2052), .CI(n1353), .CO(n1350), .S(n1351) );
  FA_X1 U896 ( .A(n2020), .B(n1355), .CI(n1358), .CO(n1352), .S(n1353) );
  HA_X1 U897 ( .A(n271), .B(n1988), .CO(n1354), .S(n1355) );
  FA_X1 U898 ( .A(n2053), .B(n1359), .CI(n2085), .CO(n1356), .S(n1357) );
  HA_X1 U899 ( .A(n2021), .B(n1362), .CO(n1358), .S(n1359) );
  FA_X1 U900 ( .A(n1363), .B(n2054), .CI(n2086), .CO(n1360), .S(n1361) );
  HA_X1 U901 ( .A(n1366), .B(n2022), .CO(n1362), .S(n1363) );
  FA_X1 U902 ( .A(n2055), .B(n1367), .CI(n1368), .CO(n1364), .S(n1365) );
  HA_X1 U903 ( .A(n2023), .B(n268), .CO(n1366), .S(n1367) );
  HA_X1 U904 ( .A(n2056), .B(n1370), .CO(n1368), .S(n1369) );
  HA_X1 U905 ( .A(n1372), .B(n2057), .CO(n1370), .S(n1371) );
  HA_X1 U906 ( .A(n265), .B(n2058), .CO(n1372), .S(n1373) );
  OAI21_X4 U907 ( .B1(n2808), .B2(n3159), .A(n2094), .ZN(n1720) );
  NAND2_X4 U908 ( .A1(n388), .A2(n484), .ZN(n2094) );
  OAI21_X4 U909 ( .B1(n2809), .B2(n3159), .A(n2095), .ZN(n717) );
  AOI21_X4 U910 ( .B1(n388), .B2(n481), .A(n1374), .ZN(n2095) );
  AND2_X4 U911 ( .A1(n333), .A2(n484), .ZN(n1374) );
  OAI21_X4 U912 ( .B1(n2810), .B2(n3159), .A(n2096), .ZN(n1721) );
  AOI222_X2 U913 ( .A1(n3149), .A2(n484), .B1(n333), .B2(n481), .C1(n388), 
        .C2(n478), .ZN(n2096) );
  OAI21_X4 U914 ( .B1(n2811), .B2(n3159), .A(n2097), .ZN(n1722) );
  AOI222_X2 U915 ( .A1(n3148), .A2(n481), .B1(n333), .B2(n478), .C1(n388), 
        .C2(n475), .ZN(n2097) );
  OAI21_X4 U916 ( .B1(n2812), .B2(n3159), .A(n2098), .ZN(n723) );
  AOI222_X2 U917 ( .A1(n3149), .A2(n478), .B1(n333), .B2(n475), .C1(n388), 
        .C2(n472), .ZN(n2098) );
  OAI21_X4 U918 ( .B1(n2813), .B2(n3159), .A(n2099), .ZN(n1723) );
  AOI222_X2 U919 ( .A1(n3148), .A2(n475), .B1(n333), .B2(n472), .C1(n388), 
        .C2(n469), .ZN(n2099) );
  OAI21_X4 U920 ( .B1(n2814), .B2(n3159), .A(n2100), .ZN(n1724) );
  AOI222_X2 U921 ( .A1(n3149), .A2(n472), .B1(n333), .B2(n469), .C1(n388), 
        .C2(n466), .ZN(n2100) );
  OAI21_X4 U922 ( .B1(n2815), .B2(n3159), .A(n2101), .ZN(n736) );
  AOI222_X2 U923 ( .A1(n3148), .A2(n469), .B1(n333), .B2(n466), .C1(n388), 
        .C2(n463), .ZN(n2101) );
  OAI21_X4 U924 ( .B1(n2816), .B2(n3159), .A(n2102), .ZN(n1725) );
  AOI222_X2 U925 ( .A1(n3149), .A2(n466), .B1(n333), .B2(n463), .C1(n388), 
        .C2(n460), .ZN(n2102) );
  OAI21_X4 U926 ( .B1(n2817), .B2(n3159), .A(n2103), .ZN(n1726) );
  AOI222_X2 U927 ( .A1(n3148), .A2(n463), .B1(n333), .B2(n460), .C1(n388), 
        .C2(n457), .ZN(n2103) );
  OAI21_X4 U928 ( .B1(n2818), .B2(n3159), .A(n2104), .ZN(n755) );
  AOI222_X2 U929 ( .A1(n3149), .A2(n460), .B1(n333), .B2(n457), .C1(n388), 
        .C2(n454), .ZN(n2104) );
  OAI21_X4 U930 ( .B1(n2819), .B2(n3159), .A(n2105), .ZN(n1727) );
  AOI222_X2 U931 ( .A1(n3148), .A2(n457), .B1(n333), .B2(n454), .C1(n388), 
        .C2(n451), .ZN(n2105) );
  OAI21_X4 U932 ( .B1(n2820), .B2(n3159), .A(n2106), .ZN(n1728) );
  AOI222_X2 U933 ( .A1(n3149), .A2(n454), .B1(n333), .B2(n451), .C1(n388), 
        .C2(n448), .ZN(n2106) );
  OAI21_X4 U934 ( .B1(n2821), .B2(n3159), .A(n2107), .ZN(n780) );
  AOI222_X2 U935 ( .A1(n3148), .A2(n451), .B1(n333), .B2(n448), .C1(n388), 
        .C2(n445), .ZN(n2107) );
  OAI21_X4 U936 ( .B1(n2822), .B2(n3159), .A(n2108), .ZN(n1729) );
  AOI222_X2 U937 ( .A1(n3149), .A2(n448), .B1(n333), .B2(n445), .C1(n388), 
        .C2(n442), .ZN(n2108) );
  OAI21_X4 U938 ( .B1(n2823), .B2(n3159), .A(n2109), .ZN(n1730) );
  AOI222_X2 U939 ( .A1(n3148), .A2(n445), .B1(n333), .B2(n442), .C1(n388), 
        .C2(n439), .ZN(n2109) );
  OAI21_X4 U940 ( .B1(n2824), .B2(n3159), .A(n2110), .ZN(n811) );
  AOI222_X2 U941 ( .A1(n3149), .A2(n442), .B1(n333), .B2(n439), .C1(n388), 
        .C2(n436), .ZN(n2110) );
  OAI21_X4 U942 ( .B1(n2825), .B2(n3159), .A(n2111), .ZN(n1731) );
  AOI222_X2 U943 ( .A1(n3149), .A2(n439), .B1(n333), .B2(n436), .C1(n388), 
        .C2(n433), .ZN(n2111) );
  OAI21_X4 U944 ( .B1(n2826), .B2(n3159), .A(n2112), .ZN(n1732) );
  AOI222_X2 U945 ( .A1(n3148), .A2(n436), .B1(n333), .B2(n433), .C1(n388), 
        .C2(n430), .ZN(n2112) );
  OAI21_X4 U946 ( .B1(n2827), .B2(n3159), .A(n2113), .ZN(n848) );
  AOI222_X2 U947 ( .A1(n3148), .A2(n433), .B1(n333), .B2(n430), .C1(n388), 
        .C2(n427), .ZN(n2113) );
  OAI21_X4 U948 ( .B1(n2828), .B2(n3159), .A(n2114), .ZN(n1733) );
  AOI222_X2 U949 ( .A1(n3149), .A2(n430), .B1(n333), .B2(n427), .C1(n388), 
        .C2(n424), .ZN(n2114) );
  OAI21_X4 U950 ( .B1(n2829), .B2(n3159), .A(n2115), .ZN(n891) );
  AOI222_X2 U951 ( .A1(n3148), .A2(n427), .B1(n333), .B2(n424), .C1(n388), 
        .C2(n421), .ZN(n2115) );
  OAI21_X4 U952 ( .B1(n2830), .B2(n3159), .A(n2116), .ZN(n1734) );
  AOI222_X2 U953 ( .A1(n3149), .A2(n424), .B1(n333), .B2(n421), .C1(n388), 
        .C2(n418), .ZN(n2116) );
  OAI21_X4 U954 ( .B1(n2831), .B2(n3159), .A(n2117), .ZN(n1735) );
  AOI222_X2 U955 ( .A1(n3149), .A2(n421), .B1(n333), .B2(n418), .C1(n388), 
        .C2(n415), .ZN(n2117) );
  OAI21_X4 U956 ( .B1(n2832), .B2(n3159), .A(n2118), .ZN(n1736) );
  AOI222_X2 U957 ( .A1(n3148), .A2(n418), .B1(n333), .B2(n415), .C1(n388), 
        .C2(n412), .ZN(n2118) );
  OAI21_X4 U958 ( .B1(n2833), .B2(n3159), .A(n2119), .ZN(n941) );
  AOI222_X2 U959 ( .A1(n3148), .A2(n415), .B1(n333), .B2(n412), .C1(n388), 
        .C2(n409), .ZN(n2119) );
  OAI21_X4 U960 ( .B1(n2834), .B2(n3158), .A(n2120), .ZN(n1737) );
  AOI222_X2 U961 ( .A1(n3148), .A2(n412), .B1(n333), .B2(n409), .C1(n388), 
        .C2(n406), .ZN(n2120) );
  OAI21_X4 U962 ( .B1(n2835), .B2(n3158), .A(n2121), .ZN(n1738) );
  AOI222_X2 U963 ( .A1(n3149), .A2(n409), .B1(n333), .B2(n406), .C1(n388), 
        .C2(n403), .ZN(n2121) );
  OAI21_X4 U964 ( .B1(n2836), .B2(n3158), .A(n2122), .ZN(n1739) );
  AOI222_X2 U965 ( .A1(n3149), .A2(n406), .B1(n333), .B2(n403), .C1(n388), 
        .C2(n400), .ZN(n2122) );
  OAI21_X4 U966 ( .B1(n2837), .B2(n3158), .A(n2123), .ZN(n1740) );
  AOI222_X2 U967 ( .A1(n3148), .A2(n403), .B1(n333), .B2(n400), .C1(n388), 
        .C2(n397), .ZN(n2123) );
  OAI21_X4 U968 ( .B1(n2838), .B2(n3158), .A(n2124), .ZN(n1741) );
  AOI222_X2 U969 ( .A1(n3149), .A2(n400), .B1(n333), .B2(n397), .C1(n388), 
        .C2(n393), .ZN(n2124) );
  OAI21_X4 U970 ( .B1(n2839), .B2(n3158), .A(n2125), .ZN(n1742) );
  AOI222_X2 U971 ( .A1(n3149), .A2(n397), .B1(n333), .B2(n393), .C1(n388), 
        .C2(n390), .ZN(n2125) );
  OAI21_X4 U972 ( .B1(n2840), .B2(n3158), .A(n2126), .ZN(n1743) );
  OAI21_X4 U974 ( .B1(n2841), .B2(n3158), .A(n2127), .ZN(n1744) );
  AND2_X4 U976 ( .A1(n3148), .A2(n390), .ZN(n1376) );
  XOR2_X2 U978 ( .A(n2128), .B(n289), .Z(n1746) );
  OAI21_X4 U979 ( .B1(n2808), .B2(n3156), .A(n2162), .ZN(n2128) );
  NAND2_X4 U980 ( .A1(n386), .A2(n484), .ZN(n2162) );
  XOR2_X2 U981 ( .A(n2129), .B(n289), .Z(n1747) );
  OAI21_X4 U982 ( .B1(n2809), .B2(n3156), .A(n2163), .ZN(n2129) );
  AOI21_X4 U983 ( .B1(n386), .B2(n481), .A(n1377), .ZN(n2163) );
  AND2_X4 U984 ( .A1(n331), .A2(n484), .ZN(n1377) );
  XOR2_X2 U985 ( .A(n2130), .B(n289), .Z(n1748) );
  OAI21_X4 U986 ( .B1(n2810), .B2(n3156), .A(n2164), .ZN(n2130) );
  AOI222_X2 U987 ( .A1(n3146), .A2(n484), .B1(n331), .B2(n481), .C1(n386), 
        .C2(n478), .ZN(n2164) );
  XOR2_X2 U988 ( .A(n2131), .B(n289), .Z(n1749) );
  OAI21_X4 U989 ( .B1(n2811), .B2(n3156), .A(n2165), .ZN(n2131) );
  AOI222_X2 U990 ( .A1(n3145), .A2(n481), .B1(n331), .B2(n478), .C1(n386), 
        .C2(n475), .ZN(n2165) );
  XOR2_X2 U991 ( .A(n2132), .B(n289), .Z(n1750) );
  OAI21_X4 U992 ( .B1(n2812), .B2(n3156), .A(n2166), .ZN(n2132) );
  AOI222_X2 U993 ( .A1(n3146), .A2(n478), .B1(n331), .B2(n475), .C1(n386), 
        .C2(n472), .ZN(n2166) );
  XOR2_X2 U994 ( .A(n2133), .B(n289), .Z(n1751) );
  OAI21_X4 U995 ( .B1(n2813), .B2(n3156), .A(n2167), .ZN(n2133) );
  AOI222_X2 U996 ( .A1(n3145), .A2(n475), .B1(n331), .B2(n472), .C1(n386), 
        .C2(n469), .ZN(n2167) );
  XOR2_X2 U997 ( .A(n2134), .B(n289), .Z(n1752) );
  OAI21_X4 U998 ( .B1(n2814), .B2(n3156), .A(n2168), .ZN(n2134) );
  AOI222_X2 U999 ( .A1(n3146), .A2(n472), .B1(n331), .B2(n469), .C1(n386), 
        .C2(n466), .ZN(n2168) );
  XOR2_X2 U1000 ( .A(n2135), .B(n289), .Z(n1753) );
  OAI21_X4 U1001 ( .B1(n2815), .B2(n3156), .A(n2169), .ZN(n2135) );
  AOI222_X2 U1002 ( .A1(n3145), .A2(n469), .B1(n331), .B2(n466), .C1(n386), 
        .C2(n463), .ZN(n2169) );
  XOR2_X2 U1003 ( .A(n2136), .B(n289), .Z(n1754) );
  OAI21_X4 U1004 ( .B1(n2816), .B2(n3156), .A(n2170), .ZN(n2136) );
  AOI222_X2 U1005 ( .A1(n3146), .A2(n466), .B1(n331), .B2(n463), .C1(n386), 
        .C2(n460), .ZN(n2170) );
  XOR2_X2 U1006 ( .A(n2137), .B(n289), .Z(n1755) );
  OAI21_X4 U1007 ( .B1(n2817), .B2(n3156), .A(n2171), .ZN(n2137) );
  AOI222_X2 U1008 ( .A1(n3145), .A2(n463), .B1(n331), .B2(n460), .C1(n386), 
        .C2(n457), .ZN(n2171) );
  XOR2_X2 U1009 ( .A(n2138), .B(n289), .Z(n1756) );
  OAI21_X4 U1010 ( .B1(n2818), .B2(n3156), .A(n2172), .ZN(n2138) );
  AOI222_X2 U1011 ( .A1(n3146), .A2(n460), .B1(n331), .B2(n457), .C1(n386), 
        .C2(n454), .ZN(n2172) );
  XOR2_X2 U1012 ( .A(n2139), .B(n289), .Z(n1757) );
  OAI21_X4 U1013 ( .B1(n2819), .B2(n3156), .A(n2173), .ZN(n2139) );
  AOI222_X2 U1014 ( .A1(n3146), .A2(n457), .B1(n331), .B2(n454), .C1(n386), 
        .C2(n451), .ZN(n2173) );
  XOR2_X2 U1015 ( .A(n2140), .B(n289), .Z(n1758) );
  OAI21_X4 U1016 ( .B1(n2820), .B2(n3156), .A(n2174), .ZN(n2140) );
  AOI222_X2 U1017 ( .A1(n3145), .A2(n454), .B1(n331), .B2(n451), .C1(n386), 
        .C2(n448), .ZN(n2174) );
  XOR2_X2 U1018 ( .A(n2141), .B(n289), .Z(n1759) );
  OAI21_X4 U1019 ( .B1(n2821), .B2(n3156), .A(n2175), .ZN(n2141) );
  AOI222_X2 U1020 ( .A1(n3145), .A2(n451), .B1(n331), .B2(n448), .C1(n386), 
        .C2(n445), .ZN(n2175) );
  XOR2_X2 U1021 ( .A(n2142), .B(n289), .Z(n1760) );
  OAI21_X4 U1022 ( .B1(n2822), .B2(n3156), .A(n2176), .ZN(n2142) );
  AOI222_X2 U1023 ( .A1(n3146), .A2(n448), .B1(n331), .B2(n445), .C1(n386), 
        .C2(n442), .ZN(n2176) );
  XOR2_X2 U1024 ( .A(n2143), .B(n289), .Z(n1761) );
  OAI21_X4 U1025 ( .B1(n2823), .B2(n3156), .A(n2177), .ZN(n2143) );
  AOI222_X2 U1026 ( .A1(n3145), .A2(n445), .B1(n331), .B2(n442), .C1(n386), 
        .C2(n439), .ZN(n2177) );
  XOR2_X2 U1027 ( .A(n2144), .B(n289), .Z(n1762) );
  OAI21_X4 U1028 ( .B1(n2824), .B2(n3156), .A(n2178), .ZN(n2144) );
  AOI222_X2 U1029 ( .A1(n3146), .A2(n442), .B1(n331), .B2(n439), .C1(n386), 
        .C2(n436), .ZN(n2178) );
  XOR2_X2 U1030 ( .A(n2145), .B(n289), .Z(n1763) );
  OAI21_X4 U1031 ( .B1(n2825), .B2(n3156), .A(n2179), .ZN(n2145) );
  AOI222_X2 U1032 ( .A1(n3145), .A2(n439), .B1(n331), .B2(n436), .C1(n386), 
        .C2(n433), .ZN(n2179) );
  XOR2_X2 U1033 ( .A(n2146), .B(n289), .Z(n1764) );
  OAI21_X4 U1034 ( .B1(n2826), .B2(n3156), .A(n2180), .ZN(n2146) );
  AOI222_X2 U1035 ( .A1(n3146), .A2(n436), .B1(n331), .B2(n433), .C1(n386), 
        .C2(n430), .ZN(n2180) );
  XOR2_X2 U1036 ( .A(n2147), .B(n289), .Z(n907) );
  OAI21_X4 U1037 ( .B1(n2827), .B2(n3156), .A(n2181), .ZN(n2147) );
  AOI222_X2 U1038 ( .A1(n3145), .A2(n433), .B1(n331), .B2(n430), .C1(n386), 
        .C2(n427), .ZN(n2181) );
  XOR2_X2 U1039 ( .A(n2148), .B(n289), .Z(n1765) );
  OAI21_X4 U1040 ( .B1(n2828), .B2(n3156), .A(n2182), .ZN(n2148) );
  AOI222_X2 U1041 ( .A1(n3146), .A2(n430), .B1(n331), .B2(n427), .C1(n386), 
        .C2(n424), .ZN(n2182) );
  XOR2_X2 U1042 ( .A(n2149), .B(n289), .Z(n1766) );
  OAI21_X4 U1043 ( .B1(n2829), .B2(n3156), .A(n2183), .ZN(n2149) );
  AOI222_X2 U1044 ( .A1(n3145), .A2(n427), .B1(n331), .B2(n424), .C1(n386), 
        .C2(n421), .ZN(n2183) );
  XOR2_X2 U1045 ( .A(n2150), .B(n289), .Z(n1767) );
  OAI21_X4 U1046 ( .B1(n2830), .B2(n3156), .A(n2184), .ZN(n2150) );
  AOI222_X2 U1047 ( .A1(n3146), .A2(n424), .B1(n331), .B2(n421), .C1(n386), 
        .C2(n418), .ZN(n2184) );
  XOR2_X2 U1048 ( .A(n2151), .B(n289), .Z(n1768) );
  OAI21_X4 U1049 ( .B1(n2831), .B2(n3156), .A(n2185), .ZN(n2151) );
  AOI222_X2 U1050 ( .A1(n3145), .A2(n421), .B1(n331), .B2(n418), .C1(n386), 
        .C2(n415), .ZN(n2185) );
  XOR2_X2 U1051 ( .A(n2152), .B(n289), .Z(n1769) );
  OAI21_X4 U1052 ( .B1(n2832), .B2(n3156), .A(n2186), .ZN(n2152) );
  AOI222_X2 U1053 ( .A1(n3146), .A2(n418), .B1(n331), .B2(n415), .C1(n386), 
        .C2(n412), .ZN(n2186) );
  XOR2_X2 U1054 ( .A(n2153), .B(n289), .Z(n1770) );
  OAI21_X4 U1055 ( .B1(n2833), .B2(n3156), .A(n2187), .ZN(n2153) );
  AOI222_X2 U1056 ( .A1(n3145), .A2(n415), .B1(n331), .B2(n412), .C1(n386), 
        .C2(n409), .ZN(n2187) );
  XOR2_X2 U1057 ( .A(n2154), .B(n289), .Z(n1771) );
  OAI21_X4 U1058 ( .B1(n2834), .B2(n3155), .A(n2188), .ZN(n2154) );
  AOI222_X2 U1059 ( .A1(n3146), .A2(n412), .B1(n331), .B2(n409), .C1(n386), 
        .C2(n406), .ZN(n2188) );
  XOR2_X2 U1060 ( .A(n2155), .B(n289), .Z(n1772) );
  OAI21_X4 U1061 ( .B1(n2835), .B2(n3155), .A(n2189), .ZN(n2155) );
  AOI222_X2 U1062 ( .A1(n3145), .A2(n409), .B1(n331), .B2(n406), .C1(n386), 
        .C2(n403), .ZN(n2189) );
  XOR2_X2 U1063 ( .A(n2156), .B(n289), .Z(n1773) );
  OAI21_X4 U1064 ( .B1(n2836), .B2(n3155), .A(n2190), .ZN(n2156) );
  AOI222_X2 U1065 ( .A1(n3146), .A2(n406), .B1(n331), .B2(n403), .C1(n386), 
        .C2(n400), .ZN(n2190) );
  XOR2_X2 U1066 ( .A(n2157), .B(n289), .Z(n1774) );
  OAI21_X4 U1067 ( .B1(n2837), .B2(n3155), .A(n2191), .ZN(n2157) );
  AOI222_X2 U1068 ( .A1(n3145), .A2(n403), .B1(n331), .B2(n400), .C1(n386), 
        .C2(n397), .ZN(n2191) );
  XOR2_X2 U1069 ( .A(n2158), .B(n289), .Z(n1775) );
  OAI21_X4 U1070 ( .B1(n2838), .B2(n3155), .A(n2192), .ZN(n2158) );
  AOI222_X2 U1071 ( .A1(n3146), .A2(n400), .B1(n331), .B2(n397), .C1(n386), 
        .C2(n393), .ZN(n2192) );
  XOR2_X2 U1072 ( .A(n2159), .B(n289), .Z(n1776) );
  OAI21_X4 U1073 ( .B1(n2839), .B2(n3155), .A(n2193), .ZN(n2159) );
  AOI222_X2 U1074 ( .A1(n3145), .A2(n397), .B1(n331), .B2(n393), .C1(n386), 
        .C2(n390), .ZN(n2193) );
  XOR2_X2 U1075 ( .A(n2160), .B(n289), .Z(n1777) );
  OAI21_X4 U1076 ( .B1(n2840), .B2(n3155), .A(n2194), .ZN(n2160) );
  XOR2_X2 U1078 ( .A(n2161), .B(n289), .Z(n1778) );
  OAI21_X4 U1079 ( .B1(n2841), .B2(n3155), .A(n2195), .ZN(n2161) );
  AND2_X4 U1081 ( .A1(n3145), .A2(n390), .ZN(n1379) );
  XOR2_X2 U1083 ( .A(n2196), .B(n286), .Z(n1780) );
  OAI21_X4 U1084 ( .B1(n2808), .B2(n3153), .A(n2230), .ZN(n2196) );
  NAND2_X4 U1085 ( .A1(n384), .A2(n484), .ZN(n2230) );
  XOR2_X2 U1086 ( .A(n2197), .B(n286), .Z(n1781) );
  OAI21_X4 U1087 ( .B1(n2809), .B2(n3153), .A(n2231), .ZN(n2197) );
  AOI21_X4 U1088 ( .B1(n384), .B2(n481), .A(n1380), .ZN(n2231) );
  AND2_X4 U1089 ( .A1(n329), .A2(n484), .ZN(n1380) );
  XOR2_X2 U1090 ( .A(n2198), .B(n286), .Z(n1782) );
  OAI21_X4 U1091 ( .B1(n2810), .B2(n3153), .A(n2232), .ZN(n2198) );
  AOI222_X2 U1092 ( .A1(n3143), .A2(n484), .B1(n329), .B2(n481), .C1(n384), 
        .C2(n478), .ZN(n2232) );
  XOR2_X2 U1093 ( .A(n2199), .B(n286), .Z(n1783) );
  OAI21_X4 U1094 ( .B1(n2811), .B2(n3153), .A(n2233), .ZN(n2199) );
  AOI222_X2 U1095 ( .A1(n3142), .A2(n481), .B1(n329), .B2(n478), .C1(n384), 
        .C2(n475), .ZN(n2233) );
  XOR2_X2 U1096 ( .A(n2200), .B(n286), .Z(n1784) );
  OAI21_X4 U1097 ( .B1(n2812), .B2(n3153), .A(n2234), .ZN(n2200) );
  AOI222_X2 U1098 ( .A1(n3143), .A2(n478), .B1(n329), .B2(n475), .C1(n384), 
        .C2(n472), .ZN(n2234) );
  XOR2_X2 U1099 ( .A(n2201), .B(n286), .Z(n1785) );
  OAI21_X4 U1100 ( .B1(n2813), .B2(n3153), .A(n2235), .ZN(n2201) );
  AOI222_X2 U1101 ( .A1(n3142), .A2(n475), .B1(n329), .B2(n472), .C1(n384), 
        .C2(n469), .ZN(n2235) );
  XOR2_X2 U1102 ( .A(n2202), .B(n286), .Z(n1786) );
  OAI21_X4 U1103 ( .B1(n2814), .B2(n3153), .A(n2236), .ZN(n2202) );
  AOI222_X2 U1104 ( .A1(n3143), .A2(n472), .B1(n329), .B2(n469), .C1(n384), 
        .C2(n466), .ZN(n2236) );
  XOR2_X2 U1105 ( .A(n2203), .B(n286), .Z(n1787) );
  OAI21_X4 U1106 ( .B1(n2815), .B2(n3153), .A(n2237), .ZN(n2203) );
  AOI222_X2 U1107 ( .A1(n3142), .A2(n469), .B1(n329), .B2(n466), .C1(n384), 
        .C2(n463), .ZN(n2237) );
  XOR2_X2 U1108 ( .A(n2204), .B(n286), .Z(n1788) );
  OAI21_X4 U1109 ( .B1(n2816), .B2(n3153), .A(n2238), .ZN(n2204) );
  AOI222_X2 U1110 ( .A1(n3143), .A2(n466), .B1(n329), .B2(n463), .C1(n384), 
        .C2(n460), .ZN(n2238) );
  XOR2_X2 U1111 ( .A(n2205), .B(n286), .Z(n1789) );
  OAI21_X4 U1112 ( .B1(n2817), .B2(n3153), .A(n2239), .ZN(n2205) );
  AOI222_X2 U1113 ( .A1(n3142), .A2(n463), .B1(n329), .B2(n460), .C1(n384), 
        .C2(n457), .ZN(n2239) );
  XOR2_X2 U1114 ( .A(n2206), .B(n286), .Z(n1790) );
  OAI21_X4 U1115 ( .B1(n2818), .B2(n3153), .A(n2240), .ZN(n2206) );
  AOI222_X2 U1116 ( .A1(n3143), .A2(n460), .B1(n329), .B2(n457), .C1(n384), 
        .C2(n454), .ZN(n2240) );
  XOR2_X2 U1117 ( .A(n2207), .B(n286), .Z(n1791) );
  OAI21_X4 U1118 ( .B1(n2819), .B2(n3153), .A(n2241), .ZN(n2207) );
  AOI222_X2 U1119 ( .A1(n3142), .A2(n457), .B1(n329), .B2(n454), .C1(n384), 
        .C2(n451), .ZN(n2241) );
  XOR2_X2 U1120 ( .A(n2208), .B(n286), .Z(n1792) );
  OAI21_X4 U1121 ( .B1(n2820), .B2(n3153), .A(n2242), .ZN(n2208) );
  AOI222_X2 U1122 ( .A1(n3143), .A2(n454), .B1(n329), .B2(n451), .C1(n384), 
        .C2(n448), .ZN(n2242) );
  XOR2_X2 U1123 ( .A(n2209), .B(n286), .Z(n1793) );
  OAI21_X4 U1124 ( .B1(n2821), .B2(n3153), .A(n2243), .ZN(n2209) );
  AOI222_X2 U1125 ( .A1(n3142), .A2(n451), .B1(n329), .B2(n448), .C1(n384), 
        .C2(n445), .ZN(n2243) );
  XOR2_X2 U1126 ( .A(n2210), .B(n286), .Z(n1794) );
  OAI21_X4 U1127 ( .B1(n2822), .B2(n3153), .A(n2244), .ZN(n2210) );
  AOI222_X2 U1128 ( .A1(n3143), .A2(n448), .B1(n329), .B2(n445), .C1(n384), 
        .C2(n442), .ZN(n2244) );
  XOR2_X2 U1129 ( .A(n2211), .B(n286), .Z(n1795) );
  OAI21_X4 U1130 ( .B1(n2823), .B2(n3153), .A(n2245), .ZN(n2211) );
  AOI222_X2 U1131 ( .A1(n3142), .A2(n445), .B1(n329), .B2(n442), .C1(n384), 
        .C2(n439), .ZN(n2245) );
  XOR2_X2 U1132 ( .A(n2212), .B(n286), .Z(n1796) );
  OAI21_X4 U1133 ( .B1(n2824), .B2(n3153), .A(n2246), .ZN(n2212) );
  AOI222_X2 U1134 ( .A1(n3143), .A2(n442), .B1(n329), .B2(n439), .C1(n384), 
        .C2(n436), .ZN(n2246) );
  XOR2_X2 U1135 ( .A(n2213), .B(n286), .Z(n1797) );
  OAI21_X4 U1136 ( .B1(n2825), .B2(n3153), .A(n2247), .ZN(n2213) );
  AOI222_X2 U1137 ( .A1(n3142), .A2(n439), .B1(n329), .B2(n436), .C1(n384), 
        .C2(n433), .ZN(n2247) );
  XOR2_X2 U1138 ( .A(n2214), .B(n286), .Z(n1798) );
  OAI21_X4 U1139 ( .B1(n2826), .B2(n3153), .A(n2248), .ZN(n2214) );
  AOI222_X2 U1140 ( .A1(n3143), .A2(n436), .B1(n329), .B2(n433), .C1(n384), 
        .C2(n430), .ZN(n2248) );
  XOR2_X2 U1141 ( .A(n2215), .B(n286), .Z(n1799) );
  OAI21_X4 U1142 ( .B1(n2827), .B2(n3153), .A(n2249), .ZN(n2215) );
  AOI222_X2 U1143 ( .A1(n3142), .A2(n433), .B1(n329), .B2(n430), .C1(n384), 
        .C2(n427), .ZN(n2249) );
  XOR2_X2 U1144 ( .A(n2216), .B(n286), .Z(n1800) );
  OAI21_X4 U1145 ( .B1(n2828), .B2(n3153), .A(n2250), .ZN(n2216) );
  AOI222_X2 U1146 ( .A1(n3143), .A2(n430), .B1(n329), .B2(n427), .C1(n384), 
        .C2(n424), .ZN(n2250) );
  XOR2_X2 U1147 ( .A(n2217), .B(n286), .Z(n1801) );
  OAI21_X4 U1148 ( .B1(n2829), .B2(n3153), .A(n2251), .ZN(n2217) );
  AOI222_X2 U1149 ( .A1(n3142), .A2(n427), .B1(n329), .B2(n424), .C1(n384), 
        .C2(n421), .ZN(n2251) );
  XOR2_X2 U1150 ( .A(n2218), .B(n286), .Z(n1802) );
  OAI21_X4 U1151 ( .B1(n2830), .B2(n3153), .A(n2252), .ZN(n2218) );
  AOI222_X2 U1152 ( .A1(n3143), .A2(n424), .B1(n329), .B2(n421), .C1(n384), 
        .C2(n418), .ZN(n2252) );
  XOR2_X2 U1153 ( .A(n2219), .B(n286), .Z(n1803) );
  OAI21_X4 U1154 ( .B1(n2831), .B2(n3153), .A(n2253), .ZN(n2219) );
  AOI222_X2 U1155 ( .A1(n3142), .A2(n421), .B1(n329), .B2(n418), .C1(n384), 
        .C2(n415), .ZN(n2253) );
  XOR2_X2 U1156 ( .A(n2220), .B(n286), .Z(n1804) );
  OAI21_X4 U1157 ( .B1(n2832), .B2(n3153), .A(n2254), .ZN(n2220) );
  AOI222_X2 U1158 ( .A1(n3143), .A2(n418), .B1(n329), .B2(n415), .C1(n384), 
        .C2(n412), .ZN(n2254) );
  XOR2_X2 U1159 ( .A(n2221), .B(n286), .Z(n1805) );
  OAI21_X4 U1160 ( .B1(n2833), .B2(n3153), .A(n2255), .ZN(n2221) );
  AOI222_X2 U1161 ( .A1(n3142), .A2(n415), .B1(n329), .B2(n412), .C1(n384), 
        .C2(n409), .ZN(n2255) );
  XOR2_X2 U1162 ( .A(n2222), .B(n286), .Z(n1806) );
  OAI21_X4 U1163 ( .B1(n2834), .B2(n3152), .A(n2256), .ZN(n2222) );
  AOI222_X2 U1164 ( .A1(n3143), .A2(n412), .B1(n329), .B2(n409), .C1(n384), 
        .C2(n406), .ZN(n2256) );
  XOR2_X2 U1165 ( .A(n2223), .B(n286), .Z(n1807) );
  OAI21_X4 U1166 ( .B1(n2835), .B2(n3152), .A(n2257), .ZN(n2223) );
  AOI222_X2 U1167 ( .A1(n3143), .A2(n409), .B1(n329), .B2(n406), .C1(n384), 
        .C2(n403), .ZN(n2257) );
  XOR2_X2 U1168 ( .A(n2224), .B(n286), .Z(n1808) );
  OAI21_X4 U1169 ( .B1(n2836), .B2(n3152), .A(n2258), .ZN(n2224) );
  AOI222_X2 U1170 ( .A1(n3142), .A2(n406), .B1(n329), .B2(n403), .C1(n384), 
        .C2(n400), .ZN(n2258) );
  XOR2_X2 U1171 ( .A(n2225), .B(n286), .Z(n1809) );
  OAI21_X4 U1172 ( .B1(n2837), .B2(n3152), .A(n2259), .ZN(n2225) );
  AOI222_X2 U1173 ( .A1(n3142), .A2(n403), .B1(n329), .B2(n400), .C1(n384), 
        .C2(n397), .ZN(n2259) );
  XOR2_X2 U1174 ( .A(n2226), .B(n286), .Z(n1810) );
  OAI21_X4 U1175 ( .B1(n2838), .B2(n3152), .A(n2260), .ZN(n2226) );
  AOI222_X2 U1176 ( .A1(n3143), .A2(n400), .B1(n329), .B2(n397), .C1(n384), 
        .C2(n393), .ZN(n2260) );
  XOR2_X2 U1177 ( .A(n2227), .B(n286), .Z(n1811) );
  OAI21_X4 U1178 ( .B1(n2839), .B2(n3152), .A(n2261), .ZN(n2227) );
  AOI222_X2 U1179 ( .A1(n3142), .A2(n397), .B1(n329), .B2(n393), .C1(n384), 
        .C2(n390), .ZN(n2261) );
  XOR2_X2 U1180 ( .A(n2228), .B(n286), .Z(n1812) );
  OAI21_X4 U1181 ( .B1(n2840), .B2(n3152), .A(n2262), .ZN(n2228) );
  XOR2_X2 U1183 ( .A(n2229), .B(n286), .Z(n1813) );
  OAI21_X4 U1184 ( .B1(n2841), .B2(n3152), .A(n2263), .ZN(n2229) );
  AND2_X4 U1186 ( .A1(n3142), .A2(n390), .ZN(n1382) );
  XOR2_X2 U1188 ( .A(n2264), .B(n283), .Z(n1815) );
  OAI21_X4 U1189 ( .B1(n2808), .B2(n3150), .A(n2298), .ZN(n2264) );
  NAND2_X4 U1190 ( .A1(n382), .A2(n484), .ZN(n2298) );
  XOR2_X2 U1191 ( .A(n2265), .B(n283), .Z(n1816) );
  OAI21_X4 U1192 ( .B1(n2809), .B2(n3150), .A(n2299), .ZN(n2265) );
  AOI21_X4 U1193 ( .B1(n382), .B2(n481), .A(n1383), .ZN(n2299) );
  AND2_X4 U1194 ( .A1(n327), .A2(n484), .ZN(n1383) );
  XOR2_X2 U1195 ( .A(n2266), .B(n283), .Z(n1817) );
  OAI21_X4 U1196 ( .B1(n2810), .B2(n357), .A(n2300), .ZN(n2266) );
  AOI222_X2 U1197 ( .A1(n3140), .A2(n484), .B1(n327), .B2(n481), .C1(n382), 
        .C2(n478), .ZN(n2300) );
  XOR2_X2 U1198 ( .A(n2267), .B(n283), .Z(n1818) );
  OAI21_X4 U1199 ( .B1(n2811), .B2(n357), .A(n2301), .ZN(n2267) );
  AOI222_X2 U1200 ( .A1(n3139), .A2(n481), .B1(n327), .B2(n478), .C1(n382), 
        .C2(n475), .ZN(n2301) );
  XOR2_X2 U1201 ( .A(n2268), .B(n283), .Z(n1819) );
  OAI21_X4 U1202 ( .B1(n2812), .B2(n357), .A(n2302), .ZN(n2268) );
  AOI222_X2 U1203 ( .A1(n3140), .A2(n478), .B1(n327), .B2(n475), .C1(n382), 
        .C2(n472), .ZN(n2302) );
  XOR2_X2 U1204 ( .A(n2269), .B(n283), .Z(n1820) );
  OAI21_X4 U1205 ( .B1(n2813), .B2(n357), .A(n2303), .ZN(n2269) );
  AOI222_X2 U1206 ( .A1(n3139), .A2(n475), .B1(n327), .B2(n472), .C1(n382), 
        .C2(n469), .ZN(n2303) );
  XOR2_X2 U1207 ( .A(n2270), .B(n283), .Z(n1821) );
  OAI21_X4 U1208 ( .B1(n2814), .B2(n357), .A(n2304), .ZN(n2270) );
  AOI222_X2 U1209 ( .A1(n3140), .A2(n472), .B1(n327), .B2(n469), .C1(n382), 
        .C2(n466), .ZN(n2304) );
  XOR2_X2 U1210 ( .A(n2271), .B(n283), .Z(n1822) );
  OAI21_X4 U1211 ( .B1(n2815), .B2(n357), .A(n2305), .ZN(n2271) );
  AOI222_X2 U1212 ( .A1(n3139), .A2(n469), .B1(n327), .B2(n466), .C1(n382), 
        .C2(n463), .ZN(n2305) );
  XOR2_X2 U1213 ( .A(n2272), .B(n283), .Z(n1823) );
  OAI21_X4 U1214 ( .B1(n2816), .B2(n357), .A(n2306), .ZN(n2272) );
  AOI222_X2 U1215 ( .A1(n3140), .A2(n466), .B1(n327), .B2(n463), .C1(n382), 
        .C2(n460), .ZN(n2306) );
  XOR2_X2 U1216 ( .A(n2273), .B(n283), .Z(n1824) );
  OAI21_X4 U1217 ( .B1(n2817), .B2(n357), .A(n2307), .ZN(n2273) );
  AOI222_X2 U1218 ( .A1(n3139), .A2(n463), .B1(n327), .B2(n460), .C1(n382), 
        .C2(n457), .ZN(n2307) );
  XOR2_X2 U1219 ( .A(n2274), .B(n283), .Z(n1825) );
  OAI21_X4 U1220 ( .B1(n2818), .B2(n357), .A(n2308), .ZN(n2274) );
  AOI222_X2 U1221 ( .A1(n3140), .A2(n460), .B1(n327), .B2(n457), .C1(n382), 
        .C2(n454), .ZN(n2308) );
  XOR2_X2 U1222 ( .A(n2275), .B(n283), .Z(n1826) );
  OAI21_X4 U1223 ( .B1(n2819), .B2(n357), .A(n2309), .ZN(n2275) );
  AOI222_X2 U1224 ( .A1(n3139), .A2(n457), .B1(n327), .B2(n454), .C1(n382), 
        .C2(n451), .ZN(n2309) );
  XOR2_X2 U1225 ( .A(n2276), .B(n283), .Z(n1827) );
  OAI21_X4 U1226 ( .B1(n2820), .B2(n357), .A(n2310), .ZN(n2276) );
  AOI222_X2 U1227 ( .A1(n3140), .A2(n454), .B1(n327), .B2(n451), .C1(n382), 
        .C2(n448), .ZN(n2310) );
  XOR2_X2 U1228 ( .A(n2277), .B(n283), .Z(n1828) );
  OAI21_X4 U1229 ( .B1(n2821), .B2(n357), .A(n2311), .ZN(n2277) );
  AOI222_X2 U1230 ( .A1(n3139), .A2(n451), .B1(n327), .B2(n448), .C1(n382), 
        .C2(n445), .ZN(n2311) );
  XOR2_X2 U1231 ( .A(n2278), .B(n283), .Z(n1829) );
  OAI21_X4 U1232 ( .B1(n2822), .B2(n357), .A(n2312), .ZN(n2278) );
  AOI222_X2 U1233 ( .A1(n3140), .A2(n448), .B1(n327), .B2(n445), .C1(n382), 
        .C2(n442), .ZN(n2312) );
  XOR2_X2 U1234 ( .A(n2279), .B(n283), .Z(n1830) );
  OAI21_X4 U1235 ( .B1(n2823), .B2(n357), .A(n2313), .ZN(n2279) );
  AOI222_X2 U1236 ( .A1(n3139), .A2(n445), .B1(n327), .B2(n442), .C1(n382), 
        .C2(n439), .ZN(n2313) );
  XOR2_X2 U1237 ( .A(n2280), .B(n283), .Z(n1831) );
  OAI21_X4 U1238 ( .B1(n2824), .B2(n357), .A(n2314), .ZN(n2280) );
  AOI222_X2 U1239 ( .A1(n3140), .A2(n442), .B1(n327), .B2(n439), .C1(n382), 
        .C2(n436), .ZN(n2314) );
  XOR2_X2 U1240 ( .A(n2281), .B(n283), .Z(n1832) );
  OAI21_X4 U1241 ( .B1(n2825), .B2(n357), .A(n2315), .ZN(n2281) );
  AOI222_X2 U1242 ( .A1(n3139), .A2(n439), .B1(n327), .B2(n436), .C1(n382), 
        .C2(n433), .ZN(n2315) );
  XOR2_X2 U1243 ( .A(n2282), .B(n283), .Z(n1833) );
  OAI21_X4 U1244 ( .B1(n2826), .B2(n357), .A(n2316), .ZN(n2282) );
  AOI222_X2 U1245 ( .A1(n3140), .A2(n436), .B1(n327), .B2(n433), .C1(n382), 
        .C2(n430), .ZN(n2316) );
  XOR2_X2 U1246 ( .A(n2283), .B(n283), .Z(n1834) );
  OAI21_X4 U1247 ( .B1(n2827), .B2(n357), .A(n2317), .ZN(n2283) );
  AOI222_X2 U1248 ( .A1(n3139), .A2(n433), .B1(n327), .B2(n430), .C1(n382), 
        .C2(n427), .ZN(n2317) );
  XOR2_X2 U1249 ( .A(n2284), .B(n283), .Z(n1835) );
  OAI21_X4 U1250 ( .B1(n2828), .B2(n357), .A(n2318), .ZN(n2284) );
  AOI222_X2 U1251 ( .A1(n3140), .A2(n430), .B1(n327), .B2(n427), .C1(n382), 
        .C2(n424), .ZN(n2318) );
  XOR2_X2 U1252 ( .A(n2285), .B(n283), .Z(n1836) );
  OAI21_X4 U1253 ( .B1(n2829), .B2(n357), .A(n2319), .ZN(n2285) );
  AOI222_X2 U1254 ( .A1(n3140), .A2(n427), .B1(n327), .B2(n424), .C1(n382), 
        .C2(n421), .ZN(n2319) );
  XOR2_X2 U1255 ( .A(n2286), .B(n283), .Z(n1837) );
  OAI21_X4 U1256 ( .B1(n2830), .B2(n357), .A(n2320), .ZN(n2286) );
  AOI222_X2 U1257 ( .A1(n3139), .A2(n424), .B1(n327), .B2(n421), .C1(n382), 
        .C2(n418), .ZN(n2320) );
  XOR2_X2 U1258 ( .A(n2287), .B(n283), .Z(n1838) );
  OAI21_X4 U1259 ( .B1(n2831), .B2(n357), .A(n2321), .ZN(n2287) );
  AOI222_X2 U1260 ( .A1(n3139), .A2(n421), .B1(n327), .B2(n418), .C1(n382), 
        .C2(n415), .ZN(n2321) );
  XOR2_X2 U1261 ( .A(n2288), .B(n283), .Z(n1839) );
  OAI21_X4 U1262 ( .B1(n2832), .B2(n357), .A(n2322), .ZN(n2288) );
  AOI222_X2 U1263 ( .A1(n3139), .A2(n418), .B1(n327), .B2(n415), .C1(n382), 
        .C2(n412), .ZN(n2322) );
  XOR2_X2 U1264 ( .A(n2289), .B(n283), .Z(n1840) );
  OAI21_X4 U1265 ( .B1(n2833), .B2(n357), .A(n2323), .ZN(n2289) );
  AOI222_X2 U1266 ( .A1(n3140), .A2(n415), .B1(n327), .B2(n412), .C1(n382), 
        .C2(n409), .ZN(n2323) );
  XOR2_X2 U1267 ( .A(n2290), .B(n283), .Z(n1841) );
  OAI21_X4 U1268 ( .B1(n2834), .B2(n357), .A(n2324), .ZN(n2290) );
  AOI222_X2 U1269 ( .A1(n3140), .A2(n412), .B1(n327), .B2(n409), .C1(n382), 
        .C2(n406), .ZN(n2324) );
  XOR2_X2 U1270 ( .A(n2291), .B(n283), .Z(n1842) );
  OAI21_X4 U1271 ( .B1(n2835), .B2(n357), .A(n2325), .ZN(n2291) );
  AOI222_X2 U1272 ( .A1(n3140), .A2(n409), .B1(n327), .B2(n406), .C1(n382), 
        .C2(n403), .ZN(n2325) );
  XOR2_X2 U1273 ( .A(n2292), .B(n283), .Z(n1843) );
  OAI21_X4 U1274 ( .B1(n2836), .B2(n357), .A(n2326), .ZN(n2292) );
  AOI222_X2 U1275 ( .A1(n3139), .A2(n406), .B1(n327), .B2(n403), .C1(n382), 
        .C2(n400), .ZN(n2326) );
  XOR2_X2 U1276 ( .A(n2293), .B(n283), .Z(n1844) );
  OAI21_X4 U1277 ( .B1(n2837), .B2(n357), .A(n2327), .ZN(n2293) );
  AOI222_X2 U1278 ( .A1(n3139), .A2(n403), .B1(n327), .B2(n400), .C1(n382), 
        .C2(n397), .ZN(n2327) );
  XOR2_X2 U1279 ( .A(n2294), .B(n283), .Z(n1845) );
  OAI21_X4 U1280 ( .B1(n2838), .B2(n357), .A(n2328), .ZN(n2294) );
  AOI222_X2 U1281 ( .A1(n3140), .A2(n400), .B1(n327), .B2(n397), .C1(n382), 
        .C2(n393), .ZN(n2328) );
  XOR2_X2 U1282 ( .A(n2295), .B(n283), .Z(n1846) );
  OAI21_X4 U1283 ( .B1(n2839), .B2(n357), .A(n2329), .ZN(n2295) );
  AOI222_X2 U1284 ( .A1(n3139), .A2(n397), .B1(n327), .B2(n393), .C1(n382), 
        .C2(n390), .ZN(n2329) );
  XOR2_X2 U1285 ( .A(n2296), .B(n283), .Z(n1847) );
  OAI21_X4 U1286 ( .B1(n2840), .B2(n357), .A(n2330), .ZN(n2296) );
  XOR2_X2 U1288 ( .A(n2297), .B(n283), .Z(n1848) );
  OAI21_X4 U1289 ( .B1(n2841), .B2(n357), .A(n2331), .ZN(n2297) );
  AND2_X4 U1291 ( .A1(n3139), .A2(n390), .ZN(n1385) );
  XOR2_X2 U1293 ( .A(n2332), .B(n280), .Z(n1850) );
  OAI21_X4 U1294 ( .B1(n2808), .B2(n3130), .A(n2366), .ZN(n2332) );
  NAND2_X4 U1295 ( .A1(n380), .A2(n484), .ZN(n2366) );
  XOR2_X2 U1296 ( .A(n2333), .B(n280), .Z(n1851) );
  OAI21_X4 U1297 ( .B1(n2809), .B2(n3130), .A(n2367), .ZN(n2333) );
  AOI21_X4 U1298 ( .B1(n380), .B2(n481), .A(n1386), .ZN(n2367) );
  AND2_X4 U1299 ( .A1(n325), .A2(n484), .ZN(n1386) );
  XOR2_X2 U1300 ( .A(n2334), .B(n280), .Z(n1852) );
  OAI21_X4 U1301 ( .B1(n2810), .B2(n354), .A(n2368), .ZN(n2334) );
  AOI222_X2 U1302 ( .A1(n3137), .A2(n484), .B1(n325), .B2(n481), .C1(n380), 
        .C2(n478), .ZN(n2368) );
  XOR2_X2 U1303 ( .A(n2335), .B(n280), .Z(n1853) );
  OAI21_X4 U1304 ( .B1(n2811), .B2(n354), .A(n2369), .ZN(n2335) );
  AOI222_X2 U1305 ( .A1(n3137), .A2(n481), .B1(n325), .B2(n478), .C1(n380), 
        .C2(n475), .ZN(n2369) );
  XOR2_X2 U1306 ( .A(n2336), .B(n280), .Z(n1854) );
  OAI21_X4 U1307 ( .B1(n2812), .B2(n354), .A(n2370), .ZN(n2336) );
  AOI222_X2 U1308 ( .A1(n3137), .A2(n478), .B1(n325), .B2(n475), .C1(n380), 
        .C2(n472), .ZN(n2370) );
  XOR2_X2 U1309 ( .A(n2337), .B(n280), .Z(n1855) );
  OAI21_X4 U1310 ( .B1(n2813), .B2(n354), .A(n2371), .ZN(n2337) );
  AOI222_X2 U1311 ( .A1(n3137), .A2(n475), .B1(n325), .B2(n472), .C1(n380), 
        .C2(n469), .ZN(n2371) );
  XOR2_X2 U1312 ( .A(n2338), .B(n280), .Z(n1856) );
  OAI21_X4 U1313 ( .B1(n2814), .B2(n354), .A(n2372), .ZN(n2338) );
  AOI222_X2 U1314 ( .A1(n3137), .A2(n472), .B1(n325), .B2(n469), .C1(n380), 
        .C2(n466), .ZN(n2372) );
  XOR2_X2 U1315 ( .A(n2339), .B(n280), .Z(n1857) );
  OAI21_X4 U1316 ( .B1(n2815), .B2(n354), .A(n2373), .ZN(n2339) );
  AOI222_X2 U1317 ( .A1(n3137), .A2(n469), .B1(n325), .B2(n466), .C1(n380), 
        .C2(n463), .ZN(n2373) );
  XOR2_X2 U1318 ( .A(n2340), .B(n280), .Z(n1858) );
  OAI21_X4 U1319 ( .B1(n2816), .B2(n354), .A(n2374), .ZN(n2340) );
  AOI222_X2 U1320 ( .A1(n3137), .A2(n466), .B1(n325), .B2(n463), .C1(n380), 
        .C2(n460), .ZN(n2374) );
  XOR2_X2 U1321 ( .A(n2341), .B(n280), .Z(n1859) );
  OAI21_X4 U1322 ( .B1(n2817), .B2(n354), .A(n2375), .ZN(n2341) );
  AOI222_X2 U1323 ( .A1(n3137), .A2(n463), .B1(n325), .B2(n460), .C1(n380), 
        .C2(n457), .ZN(n2375) );
  XOR2_X2 U1324 ( .A(n2342), .B(n280), .Z(n1860) );
  OAI21_X4 U1325 ( .B1(n2818), .B2(n354), .A(n2376), .ZN(n2342) );
  AOI222_X2 U1326 ( .A1(n3137), .A2(n460), .B1(n325), .B2(n457), .C1(n380), 
        .C2(n454), .ZN(n2376) );
  XOR2_X2 U1327 ( .A(n2343), .B(n280), .Z(n1861) );
  OAI21_X4 U1328 ( .B1(n2819), .B2(n354), .A(n2377), .ZN(n2343) );
  AOI222_X2 U1329 ( .A1(n3137), .A2(n457), .B1(n325), .B2(n454), .C1(n380), 
        .C2(n451), .ZN(n2377) );
  XOR2_X2 U1330 ( .A(n2344), .B(n280), .Z(n1862) );
  OAI21_X4 U1331 ( .B1(n2820), .B2(n354), .A(n2378), .ZN(n2344) );
  AOI222_X2 U1332 ( .A1(n3137), .A2(n454), .B1(n325), .B2(n451), .C1(n380), 
        .C2(n448), .ZN(n2378) );
  XOR2_X2 U1333 ( .A(n2345), .B(n280), .Z(n1863) );
  OAI21_X4 U1334 ( .B1(n2821), .B2(n354), .A(n2379), .ZN(n2345) );
  AOI222_X2 U1335 ( .A1(n3137), .A2(n451), .B1(n325), .B2(n448), .C1(n380), 
        .C2(n445), .ZN(n2379) );
  XOR2_X2 U1336 ( .A(n2346), .B(n280), .Z(n1864) );
  OAI21_X4 U1337 ( .B1(n2822), .B2(n354), .A(n2380), .ZN(n2346) );
  AOI222_X2 U1338 ( .A1(n3137), .A2(n448), .B1(n325), .B2(n445), .C1(n380), 
        .C2(n442), .ZN(n2380) );
  XOR2_X2 U1339 ( .A(n2347), .B(n280), .Z(n1865) );
  OAI21_X4 U1340 ( .B1(n2823), .B2(n354), .A(n2381), .ZN(n2347) );
  AOI222_X2 U1341 ( .A1(n3137), .A2(n445), .B1(n325), .B2(n442), .C1(n380), 
        .C2(n439), .ZN(n2381) );
  XOR2_X2 U1342 ( .A(n2348), .B(n280), .Z(n1866) );
  OAI21_X4 U1343 ( .B1(n2824), .B2(n354), .A(n2382), .ZN(n2348) );
  AOI222_X2 U1344 ( .A1(n3137), .A2(n442), .B1(n325), .B2(n439), .C1(n380), 
        .C2(n436), .ZN(n2382) );
  XOR2_X2 U1345 ( .A(n2349), .B(n280), .Z(n1867) );
  OAI21_X4 U1346 ( .B1(n2825), .B2(n354), .A(n2383), .ZN(n2349) );
  AOI222_X2 U1347 ( .A1(n3137), .A2(n439), .B1(n325), .B2(n436), .C1(n380), 
        .C2(n433), .ZN(n2383) );
  XOR2_X2 U1348 ( .A(n2350), .B(n280), .Z(n1868) );
  OAI21_X4 U1349 ( .B1(n2826), .B2(n354), .A(n2384), .ZN(n2350) );
  AOI222_X2 U1350 ( .A1(n3137), .A2(n436), .B1(n325), .B2(n433), .C1(n380), 
        .C2(n430), .ZN(n2384) );
  XOR2_X2 U1351 ( .A(n2351), .B(n280), .Z(n1869) );
  OAI21_X4 U1352 ( .B1(n2827), .B2(n354), .A(n2385), .ZN(n2351) );
  AOI222_X2 U1353 ( .A1(n3137), .A2(n433), .B1(n325), .B2(n430), .C1(n380), 
        .C2(n427), .ZN(n2385) );
  XOR2_X2 U1354 ( .A(n2352), .B(n280), .Z(n1870) );
  OAI21_X4 U1355 ( .B1(n2828), .B2(n354), .A(n2386), .ZN(n2352) );
  AOI222_X2 U1356 ( .A1(n3137), .A2(n430), .B1(n325), .B2(n427), .C1(n380), 
        .C2(n424), .ZN(n2386) );
  XOR2_X2 U1357 ( .A(n2353), .B(n280), .Z(n1871) );
  OAI21_X4 U1358 ( .B1(n2829), .B2(n354), .A(n2387), .ZN(n2353) );
  AOI222_X2 U1359 ( .A1(n3137), .A2(n427), .B1(n325), .B2(n424), .C1(n380), 
        .C2(n421), .ZN(n2387) );
  XOR2_X2 U1360 ( .A(n2354), .B(n280), .Z(n1872) );
  OAI21_X4 U1361 ( .B1(n2830), .B2(n354), .A(n2388), .ZN(n2354) );
  AOI222_X2 U1362 ( .A1(n3137), .A2(n424), .B1(n325), .B2(n421), .C1(n380), 
        .C2(n418), .ZN(n2388) );
  XOR2_X2 U1363 ( .A(n2355), .B(n280), .Z(n1873) );
  OAI21_X4 U1364 ( .B1(n2831), .B2(n354), .A(n2389), .ZN(n2355) );
  AOI222_X2 U1365 ( .A1(n3137), .A2(n421), .B1(n325), .B2(n418), .C1(n380), 
        .C2(n415), .ZN(n2389) );
  XOR2_X2 U1366 ( .A(n2356), .B(n280), .Z(n1874) );
  OAI21_X4 U1367 ( .B1(n2832), .B2(n354), .A(n2390), .ZN(n2356) );
  AOI222_X2 U1368 ( .A1(n3137), .A2(n418), .B1(n325), .B2(n415), .C1(n380), 
        .C2(n412), .ZN(n2390) );
  XOR2_X2 U1369 ( .A(n2357), .B(n280), .Z(n1875) );
  OAI21_X4 U1370 ( .B1(n2833), .B2(n354), .A(n2391), .ZN(n2357) );
  AOI222_X2 U1371 ( .A1(n3137), .A2(n415), .B1(n325), .B2(n412), .C1(n380), 
        .C2(n409), .ZN(n2391) );
  XOR2_X2 U1372 ( .A(n2358), .B(n280), .Z(n1876) );
  OAI21_X4 U1373 ( .B1(n2834), .B2(n354), .A(n2392), .ZN(n2358) );
  AOI222_X2 U1374 ( .A1(n3137), .A2(n412), .B1(n325), .B2(n409), .C1(n380), 
        .C2(n406), .ZN(n2392) );
  XOR2_X2 U1375 ( .A(n2359), .B(n280), .Z(n1877) );
  OAI21_X4 U1376 ( .B1(n2835), .B2(n354), .A(n2393), .ZN(n2359) );
  AOI222_X2 U1377 ( .A1(n3137), .A2(n409), .B1(n325), .B2(n406), .C1(n380), 
        .C2(n403), .ZN(n2393) );
  XOR2_X2 U1378 ( .A(n2360), .B(n280), .Z(n1878) );
  OAI21_X4 U1379 ( .B1(n2836), .B2(n354), .A(n2394), .ZN(n2360) );
  AOI222_X2 U1380 ( .A1(n3137), .A2(n406), .B1(n325), .B2(n403), .C1(n380), 
        .C2(n400), .ZN(n2394) );
  XOR2_X2 U1381 ( .A(n2361), .B(n280), .Z(n1879) );
  OAI21_X4 U1382 ( .B1(n2837), .B2(n354), .A(n2395), .ZN(n2361) );
  AOI222_X2 U1383 ( .A1(n303), .A2(n403), .B1(n325), .B2(n400), .C1(n380), 
        .C2(n397), .ZN(n2395) );
  XOR2_X2 U1384 ( .A(n2362), .B(n280), .Z(n1880) );
  OAI21_X4 U1385 ( .B1(n2838), .B2(n354), .A(n2396), .ZN(n2362) );
  AOI222_X2 U1386 ( .A1(n303), .A2(n400), .B1(n325), .B2(n397), .C1(n380), 
        .C2(n393), .ZN(n2396) );
  XOR2_X2 U1387 ( .A(n2363), .B(n280), .Z(n1881) );
  OAI21_X4 U1388 ( .B1(n2839), .B2(n354), .A(n2397), .ZN(n2363) );
  AOI222_X2 U1389 ( .A1(n303), .A2(n397), .B1(n325), .B2(n393), .C1(n380), 
        .C2(n390), .ZN(n2397) );
  XOR2_X2 U1390 ( .A(n2364), .B(n280), .Z(n1882) );
  OAI21_X4 U1391 ( .B1(n2840), .B2(n354), .A(n2398), .ZN(n2364) );
  XOR2_X2 U1393 ( .A(n2365), .B(n280), .Z(n1883) );
  OAI21_X4 U1394 ( .B1(n2841), .B2(n354), .A(n2399), .ZN(n2365) );
  AND2_X4 U1396 ( .A1(n303), .A2(n390), .ZN(n1388) );
  XOR2_X2 U1398 ( .A(n2400), .B(n277), .Z(n1885) );
  OAI21_X4 U1399 ( .B1(n2808), .B2(n3129), .A(n2434), .ZN(n2400) );
  NAND2_X4 U1400 ( .A1(n378), .A2(n484), .ZN(n2434) );
  XOR2_X2 U1401 ( .A(n2401), .B(n277), .Z(n1886) );
  OAI21_X4 U1402 ( .B1(n2809), .B2(n3129), .A(n2435), .ZN(n2401) );
  AOI21_X4 U1403 ( .B1(n378), .B2(n481), .A(n1389), .ZN(n2435) );
  AND2_X4 U1404 ( .A1(n323), .A2(n484), .ZN(n1389) );
  XOR2_X2 U1405 ( .A(n2402), .B(n277), .Z(n1887) );
  OAI21_X4 U1406 ( .B1(n2810), .B2(n351), .A(n2436), .ZN(n2402) );
  AOI222_X2 U1407 ( .A1(n3136), .A2(n484), .B1(n323), .B2(n481), .C1(n378), 
        .C2(n478), .ZN(n2436) );
  XOR2_X2 U1408 ( .A(n2403), .B(n277), .Z(n1888) );
  OAI21_X4 U1409 ( .B1(n2811), .B2(n351), .A(n2437), .ZN(n2403) );
  AOI222_X2 U1410 ( .A1(n3135), .A2(n481), .B1(n323), .B2(n478), .C1(n378), 
        .C2(n475), .ZN(n2437) );
  XOR2_X2 U1411 ( .A(n2404), .B(n277), .Z(n1889) );
  OAI21_X4 U1412 ( .B1(n2812), .B2(n351), .A(n2438), .ZN(n2404) );
  AOI222_X2 U1413 ( .A1(n3136), .A2(n478), .B1(n323), .B2(n475), .C1(n378), 
        .C2(n472), .ZN(n2438) );
  XOR2_X2 U1414 ( .A(n2405), .B(n277), .Z(n1890) );
  OAI21_X4 U1415 ( .B1(n2813), .B2(n351), .A(n2439), .ZN(n2405) );
  AOI222_X2 U1416 ( .A1(n3135), .A2(n475), .B1(n323), .B2(n472), .C1(n378), 
        .C2(n469), .ZN(n2439) );
  XOR2_X2 U1417 ( .A(n2406), .B(n277), .Z(n1891) );
  OAI21_X4 U1418 ( .B1(n2814), .B2(n351), .A(n2440), .ZN(n2406) );
  AOI222_X2 U1419 ( .A1(n3136), .A2(n472), .B1(n323), .B2(n469), .C1(n378), 
        .C2(n466), .ZN(n2440) );
  XOR2_X2 U1420 ( .A(n2407), .B(n277), .Z(n1892) );
  OAI21_X4 U1421 ( .B1(n2815), .B2(n351), .A(n2441), .ZN(n2407) );
  AOI222_X2 U1422 ( .A1(n3135), .A2(n469), .B1(n323), .B2(n466), .C1(n378), 
        .C2(n463), .ZN(n2441) );
  XOR2_X2 U1423 ( .A(n2408), .B(n277), .Z(n1893) );
  OAI21_X4 U1424 ( .B1(n2816), .B2(n351), .A(n2442), .ZN(n2408) );
  AOI222_X2 U1425 ( .A1(n3136), .A2(n466), .B1(n323), .B2(n463), .C1(n378), 
        .C2(n460), .ZN(n2442) );
  XOR2_X2 U1426 ( .A(n2409), .B(n277), .Z(n1894) );
  OAI21_X4 U1427 ( .B1(n2817), .B2(n351), .A(n2443), .ZN(n2409) );
  AOI222_X2 U1428 ( .A1(n3135), .A2(n463), .B1(n323), .B2(n460), .C1(n378), 
        .C2(n457), .ZN(n2443) );
  XOR2_X2 U1429 ( .A(n2410), .B(n277), .Z(n1895) );
  OAI21_X4 U1430 ( .B1(n2818), .B2(n351), .A(n2444), .ZN(n2410) );
  AOI222_X2 U1431 ( .A1(n3136), .A2(n460), .B1(n323), .B2(n457), .C1(n378), 
        .C2(n454), .ZN(n2444) );
  XOR2_X2 U1432 ( .A(n2411), .B(n277), .Z(n1896) );
  OAI21_X4 U1433 ( .B1(n2819), .B2(n351), .A(n2445), .ZN(n2411) );
  AOI222_X2 U1434 ( .A1(n3135), .A2(n457), .B1(n323), .B2(n454), .C1(n378), 
        .C2(n451), .ZN(n2445) );
  XOR2_X2 U1435 ( .A(n2412), .B(n277), .Z(n1897) );
  OAI21_X4 U1436 ( .B1(n2820), .B2(n351), .A(n2446), .ZN(n2412) );
  AOI222_X2 U1437 ( .A1(n3135), .A2(n454), .B1(n323), .B2(n451), .C1(n378), 
        .C2(n448), .ZN(n2446) );
  XOR2_X2 U1438 ( .A(n2413), .B(n277), .Z(n1898) );
  OAI21_X4 U1439 ( .B1(n2821), .B2(n351), .A(n2447), .ZN(n2413) );
  AOI222_X2 U1440 ( .A1(n3136), .A2(n451), .B1(n323), .B2(n448), .C1(n378), 
        .C2(n445), .ZN(n2447) );
  XOR2_X2 U1441 ( .A(n2414), .B(n277), .Z(n1899) );
  OAI21_X4 U1442 ( .B1(n2822), .B2(n351), .A(n2448), .ZN(n2414) );
  AOI222_X2 U1443 ( .A1(n3136), .A2(n448), .B1(n323), .B2(n445), .C1(n378), 
        .C2(n442), .ZN(n2448) );
  XOR2_X2 U1444 ( .A(n2415), .B(n277), .Z(n1900) );
  OAI21_X4 U1445 ( .B1(n2823), .B2(n351), .A(n2449), .ZN(n2415) );
  AOI222_X2 U1446 ( .A1(n3136), .A2(n445), .B1(n323), .B2(n442), .C1(n378), 
        .C2(n439), .ZN(n2449) );
  XOR2_X2 U1447 ( .A(n2416), .B(n277), .Z(n1901) );
  OAI21_X4 U1448 ( .B1(n2824), .B2(n351), .A(n2450), .ZN(n2416) );
  AOI222_X2 U1449 ( .A1(n3135), .A2(n442), .B1(n323), .B2(n439), .C1(n378), 
        .C2(n436), .ZN(n2450) );
  XOR2_X2 U1450 ( .A(n2417), .B(n277), .Z(n1902) );
  OAI21_X4 U1451 ( .B1(n2825), .B2(n351), .A(n2451), .ZN(n2417) );
  AOI222_X2 U1452 ( .A1(n3136), .A2(n439), .B1(n323), .B2(n436), .C1(n378), 
        .C2(n433), .ZN(n2451) );
  XOR2_X2 U1453 ( .A(n2418), .B(n277), .Z(n1903) );
  OAI21_X4 U1454 ( .B1(n2826), .B2(n351), .A(n2452), .ZN(n2418) );
  AOI222_X2 U1455 ( .A1(n3135), .A2(n436), .B1(n323), .B2(n433), .C1(n378), 
        .C2(n430), .ZN(n2452) );
  XOR2_X2 U1456 ( .A(n2419), .B(n277), .Z(n1904) );
  OAI21_X4 U1457 ( .B1(n2827), .B2(n351), .A(n2453), .ZN(n2419) );
  AOI222_X2 U1458 ( .A1(n3135), .A2(n433), .B1(n323), .B2(n430), .C1(n378), 
        .C2(n427), .ZN(n2453) );
  XOR2_X2 U1459 ( .A(n2420), .B(n277), .Z(n1905) );
  OAI21_X4 U1460 ( .B1(n2828), .B2(n351), .A(n2454), .ZN(n2420) );
  AOI222_X2 U1461 ( .A1(n3136), .A2(n430), .B1(n323), .B2(n427), .C1(n378), 
        .C2(n424), .ZN(n2454) );
  XOR2_X2 U1462 ( .A(n2421), .B(n277), .Z(n1906) );
  OAI21_X4 U1463 ( .B1(n2829), .B2(n351), .A(n2455), .ZN(n2421) );
  AOI222_X2 U1464 ( .A1(n3135), .A2(n427), .B1(n323), .B2(n424), .C1(n378), 
        .C2(n421), .ZN(n2455) );
  XOR2_X2 U1465 ( .A(n2422), .B(n277), .Z(n1907) );
  OAI21_X4 U1466 ( .B1(n2830), .B2(n351), .A(n2456), .ZN(n2422) );
  AOI222_X2 U1467 ( .A1(n3135), .A2(n424), .B1(n323), .B2(n421), .C1(n378), 
        .C2(n418), .ZN(n2456) );
  XOR2_X2 U1468 ( .A(n2423), .B(n277), .Z(n1908) );
  OAI21_X4 U1469 ( .B1(n2831), .B2(n351), .A(n2457), .ZN(n2423) );
  AOI222_X2 U1470 ( .A1(n3136), .A2(n421), .B1(n323), .B2(n418), .C1(n378), 
        .C2(n415), .ZN(n2457) );
  XOR2_X2 U1471 ( .A(n2424), .B(n277), .Z(n1909) );
  OAI21_X4 U1472 ( .B1(n2832), .B2(n351), .A(n2458), .ZN(n2424) );
  AOI222_X2 U1473 ( .A1(n3135), .A2(n418), .B1(n323), .B2(n415), .C1(n378), 
        .C2(n412), .ZN(n2458) );
  XOR2_X2 U1474 ( .A(n2425), .B(n277), .Z(n1910) );
  OAI21_X4 U1475 ( .B1(n2833), .B2(n351), .A(n2459), .ZN(n2425) );
  AOI222_X2 U1476 ( .A1(n3136), .A2(n415), .B1(n323), .B2(n412), .C1(n378), 
        .C2(n409), .ZN(n2459) );
  XOR2_X2 U1477 ( .A(n2426), .B(n277), .Z(n1911) );
  OAI21_X4 U1478 ( .B1(n2834), .B2(n351), .A(n2460), .ZN(n2426) );
  AOI222_X2 U1479 ( .A1(n3136), .A2(n412), .B1(n323), .B2(n409), .C1(n378), 
        .C2(n406), .ZN(n2460) );
  XOR2_X2 U1480 ( .A(n2427), .B(n277), .Z(n1912) );
  OAI21_X4 U1481 ( .B1(n2835), .B2(n351), .A(n2461), .ZN(n2427) );
  AOI222_X2 U1482 ( .A1(n3135), .A2(n409), .B1(n323), .B2(n406), .C1(n378), 
        .C2(n403), .ZN(n2461) );
  XOR2_X2 U1483 ( .A(n2428), .B(n277), .Z(n1913) );
  OAI21_X4 U1484 ( .B1(n2836), .B2(n351), .A(n2462), .ZN(n2428) );
  AOI222_X2 U1485 ( .A1(n3136), .A2(n406), .B1(n323), .B2(n403), .C1(n378), 
        .C2(n400), .ZN(n2462) );
  XOR2_X2 U1486 ( .A(n2429), .B(n277), .Z(n1914) );
  OAI21_X4 U1487 ( .B1(n2837), .B2(n351), .A(n2463), .ZN(n2429) );
  AOI222_X2 U1488 ( .A1(n3135), .A2(n403), .B1(n323), .B2(n400), .C1(n378), 
        .C2(n397), .ZN(n2463) );
  XOR2_X2 U1489 ( .A(n2430), .B(n277), .Z(n1915) );
  OAI21_X4 U1490 ( .B1(n2838), .B2(n351), .A(n2464), .ZN(n2430) );
  AOI222_X2 U1491 ( .A1(n3136), .A2(n400), .B1(n323), .B2(n397), .C1(n378), 
        .C2(n393), .ZN(n2464) );
  XOR2_X2 U1492 ( .A(n2431), .B(n277), .Z(n1916) );
  OAI21_X4 U1493 ( .B1(n2839), .B2(n351), .A(n2465), .ZN(n2431) );
  AOI222_X2 U1494 ( .A1(n3135), .A2(n397), .B1(n323), .B2(n393), .C1(n378), 
        .C2(n390), .ZN(n2465) );
  XOR2_X2 U1495 ( .A(n2432), .B(n277), .Z(n1917) );
  OAI21_X4 U1496 ( .B1(n2840), .B2(n351), .A(n2466), .ZN(n2432) );
  XOR2_X2 U1498 ( .A(n2433), .B(n277), .Z(n1918) );
  OAI21_X4 U1499 ( .B1(n2841), .B2(n351), .A(n2467), .ZN(n2433) );
  AND2_X4 U1501 ( .A1(n3135), .A2(n390), .ZN(n1391) );
  XOR2_X2 U1503 ( .A(n2468), .B(n274), .Z(n1920) );
  OAI21_X4 U1504 ( .B1(n2808), .B2(n3128), .A(n2502), .ZN(n2468) );
  NAND2_X4 U1505 ( .A1(n376), .A2(n484), .ZN(n2502) );
  XOR2_X2 U1506 ( .A(n2469), .B(n274), .Z(n1921) );
  OAI21_X4 U1507 ( .B1(n2809), .B2(n3128), .A(n2503), .ZN(n2469) );
  AOI21_X4 U1508 ( .B1(n376), .B2(n481), .A(n1392), .ZN(n2503) );
  AND2_X4 U1509 ( .A1(n321), .A2(n484), .ZN(n1392) );
  XOR2_X2 U1510 ( .A(n2470), .B(n274), .Z(n1922) );
  OAI21_X4 U1511 ( .B1(n2810), .B2(n348), .A(n2504), .ZN(n2470) );
  AOI222_X2 U1512 ( .A1(n3133), .A2(n484), .B1(n321), .B2(n481), .C1(n376), 
        .C2(n478), .ZN(n2504) );
  XOR2_X2 U1513 ( .A(n2471), .B(n274), .Z(n1923) );
  OAI21_X4 U1514 ( .B1(n2811), .B2(n348), .A(n2505), .ZN(n2471) );
  AOI222_X2 U1515 ( .A1(n3132), .A2(n481), .B1(n321), .B2(n478), .C1(n376), 
        .C2(n475), .ZN(n2505) );
  XOR2_X2 U1516 ( .A(n2472), .B(n274), .Z(n1924) );
  OAI21_X4 U1517 ( .B1(n2812), .B2(n348), .A(n2506), .ZN(n2472) );
  AOI222_X2 U1518 ( .A1(n3133), .A2(n478), .B1(n321), .B2(n475), .C1(n376), 
        .C2(n472), .ZN(n2506) );
  XOR2_X2 U1519 ( .A(n2473), .B(n274), .Z(n1925) );
  OAI21_X4 U1520 ( .B1(n2813), .B2(n348), .A(n2507), .ZN(n2473) );
  AOI222_X2 U1521 ( .A1(n3132), .A2(n475), .B1(n321), .B2(n472), .C1(n376), 
        .C2(n469), .ZN(n2507) );
  XOR2_X2 U1522 ( .A(n2474), .B(n274), .Z(n1926) );
  OAI21_X4 U1523 ( .B1(n2814), .B2(n348), .A(n2508), .ZN(n2474) );
  AOI222_X2 U1524 ( .A1(n3133), .A2(n472), .B1(n321), .B2(n469), .C1(n376), 
        .C2(n466), .ZN(n2508) );
  XOR2_X2 U1525 ( .A(n2475), .B(n274), .Z(n1927) );
  OAI21_X4 U1526 ( .B1(n2815), .B2(n348), .A(n2509), .ZN(n2475) );
  AOI222_X2 U1527 ( .A1(n3132), .A2(n469), .B1(n321), .B2(n466), .C1(n376), 
        .C2(n463), .ZN(n2509) );
  XOR2_X2 U1528 ( .A(n2476), .B(n274), .Z(n1928) );
  OAI21_X4 U1529 ( .B1(n2816), .B2(n348), .A(n2510), .ZN(n2476) );
  AOI222_X2 U1530 ( .A1(n3133), .A2(n466), .B1(n321), .B2(n463), .C1(n376), 
        .C2(n460), .ZN(n2510) );
  XOR2_X2 U1531 ( .A(n2477), .B(n274), .Z(n1929) );
  OAI21_X4 U1532 ( .B1(n2817), .B2(n348), .A(n2511), .ZN(n2477) );
  AOI222_X2 U1533 ( .A1(n3132), .A2(n463), .B1(n321), .B2(n460), .C1(n376), 
        .C2(n457), .ZN(n2511) );
  XOR2_X2 U1534 ( .A(n2478), .B(n274), .Z(n1930) );
  OAI21_X4 U1535 ( .B1(n2818), .B2(n348), .A(n2512), .ZN(n2478) );
  AOI222_X2 U1536 ( .A1(n3132), .A2(n460), .B1(n321), .B2(n457), .C1(n376), 
        .C2(n454), .ZN(n2512) );
  XOR2_X2 U1537 ( .A(n2479), .B(n274), .Z(n1931) );
  OAI21_X4 U1538 ( .B1(n2819), .B2(n348), .A(n2513), .ZN(n2479) );
  AOI222_X2 U1539 ( .A1(n3133), .A2(n457), .B1(n321), .B2(n454), .C1(n376), 
        .C2(n451), .ZN(n2513) );
  XOR2_X2 U1540 ( .A(n2480), .B(n274), .Z(n1932) );
  OAI21_X4 U1541 ( .B1(n2820), .B2(n348), .A(n2514), .ZN(n2480) );
  AOI222_X2 U1542 ( .A1(n3133), .A2(n454), .B1(n321), .B2(n451), .C1(n376), 
        .C2(n448), .ZN(n2514) );
  XOR2_X2 U1543 ( .A(n2481), .B(n274), .Z(n1933) );
  OAI21_X4 U1544 ( .B1(n2821), .B2(n348), .A(n2515), .ZN(n2481) );
  AOI222_X2 U1545 ( .A1(n3132), .A2(n451), .B1(n321), .B2(n448), .C1(n376), 
        .C2(n445), .ZN(n2515) );
  XOR2_X2 U1546 ( .A(n2482), .B(n274), .Z(n1934) );
  OAI21_X4 U1547 ( .B1(n2822), .B2(n348), .A(n2516), .ZN(n2482) );
  AOI222_X2 U1548 ( .A1(n3133), .A2(n448), .B1(n321), .B2(n445), .C1(n376), 
        .C2(n442), .ZN(n2516) );
  XOR2_X2 U1549 ( .A(n2483), .B(n274), .Z(n1935) );
  OAI21_X4 U1550 ( .B1(n2823), .B2(n348), .A(n2517), .ZN(n2483) );
  AOI222_X2 U1551 ( .A1(n3132), .A2(n445), .B1(n321), .B2(n442), .C1(n376), 
        .C2(n439), .ZN(n2517) );
  XOR2_X2 U1552 ( .A(n2484), .B(n274), .Z(n1936) );
  OAI21_X4 U1553 ( .B1(n2824), .B2(n348), .A(n2518), .ZN(n2484) );
  AOI222_X2 U1554 ( .A1(n3133), .A2(n442), .B1(n321), .B2(n439), .C1(n376), 
        .C2(n436), .ZN(n2518) );
  XOR2_X2 U1555 ( .A(n2485), .B(n274), .Z(n1937) );
  OAI21_X4 U1556 ( .B1(n2825), .B2(n348), .A(n2519), .ZN(n2485) );
  AOI222_X2 U1557 ( .A1(n3133), .A2(n439), .B1(n321), .B2(n436), .C1(n376), 
        .C2(n433), .ZN(n2519) );
  XOR2_X2 U1558 ( .A(n2486), .B(n274), .Z(n1938) );
  OAI21_X4 U1559 ( .B1(n2826), .B2(n348), .A(n2520), .ZN(n2486) );
  AOI222_X2 U1560 ( .A1(n3132), .A2(n436), .B1(n321), .B2(n433), .C1(n376), 
        .C2(n430), .ZN(n2520) );
  XOR2_X2 U1561 ( .A(n2487), .B(n274), .Z(n1939) );
  OAI21_X4 U1562 ( .B1(n2827), .B2(n348), .A(n2521), .ZN(n2487) );
  AOI222_X2 U1563 ( .A1(n3133), .A2(n433), .B1(n321), .B2(n430), .C1(n376), 
        .C2(n427), .ZN(n2521) );
  XOR2_X2 U1564 ( .A(n2488), .B(n274), .Z(n1940) );
  OAI21_X4 U1565 ( .B1(n2828), .B2(n348), .A(n2522), .ZN(n2488) );
  AOI222_X2 U1566 ( .A1(n3132), .A2(n430), .B1(n321), .B2(n427), .C1(n376), 
        .C2(n424), .ZN(n2522) );
  XOR2_X2 U1567 ( .A(n2489), .B(n274), .Z(n1941) );
  OAI21_X4 U1568 ( .B1(n2829), .B2(n348), .A(n2523), .ZN(n2489) );
  AOI222_X2 U1569 ( .A1(n3133), .A2(n427), .B1(n321), .B2(n424), .C1(n376), 
        .C2(n421), .ZN(n2523) );
  XOR2_X2 U1570 ( .A(n2490), .B(n274), .Z(n1942) );
  OAI21_X4 U1571 ( .B1(n2830), .B2(n348), .A(n2524), .ZN(n2490) );
  AOI222_X2 U1572 ( .A1(n3132), .A2(n424), .B1(n321), .B2(n421), .C1(n376), 
        .C2(n418), .ZN(n2524) );
  XOR2_X2 U1573 ( .A(n2491), .B(n274), .Z(n1943) );
  OAI21_X4 U1574 ( .B1(n2831), .B2(n348), .A(n2525), .ZN(n2491) );
  AOI222_X2 U1575 ( .A1(n3133), .A2(n421), .B1(n321), .B2(n418), .C1(n376), 
        .C2(n415), .ZN(n2525) );
  XOR2_X2 U1576 ( .A(n2492), .B(n274), .Z(n1944) );
  OAI21_X4 U1577 ( .B1(n2832), .B2(n348), .A(n2526), .ZN(n2492) );
  AOI222_X2 U1578 ( .A1(n3132), .A2(n418), .B1(n321), .B2(n415), .C1(n376), 
        .C2(n412), .ZN(n2526) );
  XOR2_X2 U1579 ( .A(n2493), .B(n274), .Z(n1945) );
  OAI21_X4 U1580 ( .B1(n2833), .B2(n348), .A(n2527), .ZN(n2493) );
  AOI222_X2 U1581 ( .A1(n3132), .A2(n415), .B1(n321), .B2(n412), .C1(n376), 
        .C2(n409), .ZN(n2527) );
  XOR2_X2 U1582 ( .A(n2494), .B(n274), .Z(n1946) );
  OAI21_X4 U1583 ( .B1(n2834), .B2(n348), .A(n2528), .ZN(n2494) );
  AOI222_X2 U1584 ( .A1(n3133), .A2(n412), .B1(n321), .B2(n409), .C1(n376), 
        .C2(n406), .ZN(n2528) );
  XOR2_X2 U1585 ( .A(n2495), .B(n274), .Z(n1947) );
  OAI21_X4 U1586 ( .B1(n2835), .B2(n348), .A(n2529), .ZN(n2495) );
  AOI222_X2 U1587 ( .A1(n3132), .A2(n409), .B1(n321), .B2(n406), .C1(n376), 
        .C2(n403), .ZN(n2529) );
  XOR2_X2 U1588 ( .A(n2496), .B(n274), .Z(n1948) );
  OAI21_X4 U1589 ( .B1(n2836), .B2(n348), .A(n2530), .ZN(n2496) );
  AOI222_X2 U1590 ( .A1(n3133), .A2(n406), .B1(n321), .B2(n403), .C1(n376), 
        .C2(n400), .ZN(n2530) );
  XOR2_X2 U1591 ( .A(n2497), .B(n274), .Z(n1949) );
  OAI21_X4 U1592 ( .B1(n2837), .B2(n348), .A(n2531), .ZN(n2497) );
  AOI222_X2 U1593 ( .A1(n3132), .A2(n403), .B1(n321), .B2(n400), .C1(n376), 
        .C2(n397), .ZN(n2531) );
  XOR2_X2 U1594 ( .A(n2498), .B(n274), .Z(n1950) );
  OAI21_X4 U1595 ( .B1(n2838), .B2(n348), .A(n2532), .ZN(n2498) );
  AOI222_X2 U1596 ( .A1(n3133), .A2(n400), .B1(n321), .B2(n397), .C1(n376), 
        .C2(n393), .ZN(n2532) );
  XOR2_X2 U1597 ( .A(n2499), .B(n274), .Z(n1951) );
  OAI21_X4 U1598 ( .B1(n2839), .B2(n348), .A(n2533), .ZN(n2499) );
  AOI222_X2 U1599 ( .A1(n3132), .A2(n397), .B1(n321), .B2(n393), .C1(n376), 
        .C2(n390), .ZN(n2533) );
  XOR2_X2 U1600 ( .A(n2500), .B(n274), .Z(n1952) );
  OAI21_X4 U1601 ( .B1(n2840), .B2(n348), .A(n2534), .ZN(n2500) );
  OAI21_X4 U1604 ( .B1(n2841), .B2(n348), .A(n2535), .ZN(n2501) );
  AND2_X4 U1606 ( .A1(n3132), .A2(n390), .ZN(n1394) );
  XOR2_X2 U1608 ( .A(n2536), .B(n271), .Z(n1955) );
  OAI21_X4 U1609 ( .B1(n2808), .B2(n345), .A(n2570), .ZN(n2536) );
  NAND2_X4 U1610 ( .A1(n374), .A2(n484), .ZN(n2570) );
  XOR2_X2 U1611 ( .A(n2537), .B(n271), .Z(n1956) );
  OAI21_X4 U1612 ( .B1(n2809), .B2(n345), .A(n2571), .ZN(n2537) );
  AOI21_X4 U1613 ( .B1(n374), .B2(n481), .A(n1395), .ZN(n2571) );
  AND2_X4 U1614 ( .A1(n319), .A2(n484), .ZN(n1395) );
  XOR2_X2 U1615 ( .A(n2538), .B(n271), .Z(n1957) );
  OAI21_X4 U1616 ( .B1(n2810), .B2(n345), .A(n2572), .ZN(n2538) );
  AOI222_X2 U1617 ( .A1(n297), .A2(n484), .B1(n319), .B2(n481), .C1(n374), 
        .C2(n478), .ZN(n2572) );
  XOR2_X2 U1618 ( .A(n2539), .B(n271), .Z(n1958) );
  OAI21_X4 U1619 ( .B1(n2811), .B2(n345), .A(n2573), .ZN(n2539) );
  AOI222_X2 U1620 ( .A1(n297), .A2(n481), .B1(n319), .B2(n478), .C1(n374), 
        .C2(n475), .ZN(n2573) );
  XOR2_X2 U1621 ( .A(n2540), .B(n271), .Z(n1959) );
  OAI21_X4 U1622 ( .B1(n2812), .B2(n345), .A(n2574), .ZN(n2540) );
  AOI222_X2 U1623 ( .A1(n297), .A2(n478), .B1(n319), .B2(n475), .C1(n374), 
        .C2(n472), .ZN(n2574) );
  XOR2_X2 U1624 ( .A(n2541), .B(n271), .Z(n1960) );
  OAI21_X4 U1625 ( .B1(n2813), .B2(n345), .A(n2575), .ZN(n2541) );
  AOI222_X2 U1626 ( .A1(n297), .A2(n475), .B1(n319), .B2(n472), .C1(n374), 
        .C2(n469), .ZN(n2575) );
  XOR2_X2 U1627 ( .A(n2542), .B(n271), .Z(n1961) );
  OAI21_X4 U1628 ( .B1(n2814), .B2(n345), .A(n2576), .ZN(n2542) );
  AOI222_X2 U1629 ( .A1(n297), .A2(n472), .B1(n319), .B2(n469), .C1(n374), 
        .C2(n466), .ZN(n2576) );
  XOR2_X2 U1630 ( .A(n2543), .B(n271), .Z(n1962) );
  OAI21_X4 U1631 ( .B1(n2815), .B2(n345), .A(n2577), .ZN(n2543) );
  AOI222_X2 U1632 ( .A1(n297), .A2(n469), .B1(n319), .B2(n466), .C1(n374), 
        .C2(n463), .ZN(n2577) );
  XOR2_X2 U1633 ( .A(n2544), .B(n271), .Z(n1963) );
  OAI21_X4 U1634 ( .B1(n2816), .B2(n345), .A(n2578), .ZN(n2544) );
  AOI222_X2 U1635 ( .A1(n297), .A2(n466), .B1(n319), .B2(n463), .C1(n374), 
        .C2(n460), .ZN(n2578) );
  XOR2_X2 U1636 ( .A(n2545), .B(n271), .Z(n1964) );
  OAI21_X4 U1637 ( .B1(n2817), .B2(n345), .A(n2579), .ZN(n2545) );
  AOI222_X2 U1638 ( .A1(n297), .A2(n463), .B1(n319), .B2(n460), .C1(n374), 
        .C2(n457), .ZN(n2579) );
  XOR2_X2 U1639 ( .A(n2546), .B(n271), .Z(n1965) );
  OAI21_X4 U1640 ( .B1(n2818), .B2(n345), .A(n2580), .ZN(n2546) );
  AOI222_X2 U1641 ( .A1(n297), .A2(n460), .B1(n319), .B2(n457), .C1(n374), 
        .C2(n454), .ZN(n2580) );
  XOR2_X2 U1642 ( .A(n2547), .B(n271), .Z(n1966) );
  OAI21_X4 U1643 ( .B1(n2819), .B2(n345), .A(n2581), .ZN(n2547) );
  AOI222_X2 U1644 ( .A1(n297), .A2(n457), .B1(n319), .B2(n454), .C1(n374), 
        .C2(n451), .ZN(n2581) );
  XOR2_X2 U1645 ( .A(n2548), .B(n271), .Z(n1967) );
  OAI21_X4 U1646 ( .B1(n2820), .B2(n345), .A(n2582), .ZN(n2548) );
  AOI222_X2 U1647 ( .A1(n297), .A2(n454), .B1(n319), .B2(n451), .C1(n374), 
        .C2(n448), .ZN(n2582) );
  XOR2_X2 U1648 ( .A(n2549), .B(n271), .Z(n1968) );
  OAI21_X4 U1649 ( .B1(n2821), .B2(n345), .A(n2583), .ZN(n2549) );
  AOI222_X2 U1650 ( .A1(n297), .A2(n451), .B1(n319), .B2(n448), .C1(n374), 
        .C2(n445), .ZN(n2583) );
  XOR2_X2 U1651 ( .A(n2550), .B(n271), .Z(n1969) );
  OAI21_X4 U1652 ( .B1(n2822), .B2(n345), .A(n2584), .ZN(n2550) );
  AOI222_X2 U1653 ( .A1(n297), .A2(n448), .B1(n319), .B2(n445), .C1(n374), 
        .C2(n442), .ZN(n2584) );
  XOR2_X2 U1654 ( .A(n2551), .B(n271), .Z(n1970) );
  OAI21_X4 U1655 ( .B1(n2823), .B2(n345), .A(n2585), .ZN(n2551) );
  AOI222_X2 U1656 ( .A1(n297), .A2(n445), .B1(n319), .B2(n442), .C1(n374), 
        .C2(n439), .ZN(n2585) );
  XOR2_X2 U1657 ( .A(n2552), .B(n271), .Z(n1971) );
  OAI21_X4 U1658 ( .B1(n2824), .B2(n345), .A(n2586), .ZN(n2552) );
  AOI222_X2 U1659 ( .A1(n297), .A2(n442), .B1(n319), .B2(n439), .C1(n374), 
        .C2(n436), .ZN(n2586) );
  XOR2_X2 U1660 ( .A(n2553), .B(n271), .Z(n1972) );
  OAI21_X4 U1661 ( .B1(n2825), .B2(n345), .A(n2587), .ZN(n2553) );
  AOI222_X2 U1662 ( .A1(n297), .A2(n439), .B1(n319), .B2(n436), .C1(n374), 
        .C2(n433), .ZN(n2587) );
  XOR2_X2 U1663 ( .A(n2554), .B(n271), .Z(n1973) );
  OAI21_X4 U1664 ( .B1(n2826), .B2(n345), .A(n2588), .ZN(n2554) );
  AOI222_X2 U1665 ( .A1(n297), .A2(n436), .B1(n319), .B2(n433), .C1(n374), 
        .C2(n430), .ZN(n2588) );
  XOR2_X2 U1666 ( .A(n2555), .B(n271), .Z(n1974) );
  OAI21_X4 U1667 ( .B1(n2827), .B2(n345), .A(n2589), .ZN(n2555) );
  AOI222_X2 U1668 ( .A1(n297), .A2(n433), .B1(n319), .B2(n430), .C1(n374), 
        .C2(n427), .ZN(n2589) );
  XOR2_X2 U1669 ( .A(n2556), .B(n271), .Z(n1975) );
  OAI21_X4 U1670 ( .B1(n2828), .B2(n345), .A(n2590), .ZN(n2556) );
  AOI222_X2 U1671 ( .A1(n297), .A2(n430), .B1(n319), .B2(n427), .C1(n374), 
        .C2(n424), .ZN(n2590) );
  XOR2_X2 U1672 ( .A(n2557), .B(n271), .Z(n1976) );
  OAI21_X4 U1673 ( .B1(n2829), .B2(n345), .A(n2591), .ZN(n2557) );
  AOI222_X2 U1674 ( .A1(n297), .A2(n427), .B1(n319), .B2(n424), .C1(n374), 
        .C2(n421), .ZN(n2591) );
  XOR2_X2 U1675 ( .A(n2558), .B(n271), .Z(n1977) );
  OAI21_X4 U1676 ( .B1(n2830), .B2(n345), .A(n2592), .ZN(n2558) );
  AOI222_X2 U1677 ( .A1(n297), .A2(n424), .B1(n319), .B2(n421), .C1(n374), 
        .C2(n418), .ZN(n2592) );
  XOR2_X2 U1678 ( .A(n2559), .B(n271), .Z(n1978) );
  OAI21_X4 U1679 ( .B1(n2831), .B2(n345), .A(n2593), .ZN(n2559) );
  AOI222_X2 U1680 ( .A1(n297), .A2(n421), .B1(n319), .B2(n418), .C1(n374), 
        .C2(n415), .ZN(n2593) );
  XOR2_X2 U1681 ( .A(n2560), .B(n271), .Z(n1979) );
  OAI21_X4 U1682 ( .B1(n2832), .B2(n345), .A(n2594), .ZN(n2560) );
  AOI222_X2 U1683 ( .A1(n297), .A2(n418), .B1(n319), .B2(n415), .C1(n374), 
        .C2(n412), .ZN(n2594) );
  XOR2_X2 U1684 ( .A(n2561), .B(n271), .Z(n1980) );
  OAI21_X4 U1685 ( .B1(n2833), .B2(n345), .A(n2595), .ZN(n2561) );
  AOI222_X2 U1686 ( .A1(n297), .A2(n415), .B1(n319), .B2(n412), .C1(n374), 
        .C2(n409), .ZN(n2595) );
  XOR2_X2 U1687 ( .A(n2562), .B(n271), .Z(n1981) );
  OAI21_X4 U1688 ( .B1(n2834), .B2(n345), .A(n2596), .ZN(n2562) );
  AOI222_X2 U1689 ( .A1(n297), .A2(n412), .B1(n319), .B2(n409), .C1(n374), 
        .C2(n406), .ZN(n2596) );
  XOR2_X2 U1690 ( .A(n2563), .B(n271), .Z(n1982) );
  OAI21_X4 U1691 ( .B1(n2835), .B2(n345), .A(n2597), .ZN(n2563) );
  AOI222_X2 U1692 ( .A1(n297), .A2(n409), .B1(n319), .B2(n406), .C1(n374), 
        .C2(n403), .ZN(n2597) );
  XOR2_X2 U1693 ( .A(n2564), .B(n271), .Z(n1983) );
  OAI21_X4 U1694 ( .B1(n2836), .B2(n345), .A(n2598), .ZN(n2564) );
  AOI222_X2 U1695 ( .A1(n297), .A2(n406), .B1(n319), .B2(n403), .C1(n374), 
        .C2(n400), .ZN(n2598) );
  XOR2_X2 U1696 ( .A(n2565), .B(n271), .Z(n1984) );
  OAI21_X4 U1697 ( .B1(n2837), .B2(n345), .A(n2599), .ZN(n2565) );
  AOI222_X2 U1698 ( .A1(n297), .A2(n403), .B1(n319), .B2(n400), .C1(n374), 
        .C2(n397), .ZN(n2599) );
  XOR2_X2 U1699 ( .A(n2566), .B(n271), .Z(n1985) );
  OAI21_X4 U1700 ( .B1(n2838), .B2(n345), .A(n2600), .ZN(n2566) );
  AOI222_X2 U1701 ( .A1(n297), .A2(n400), .B1(n319), .B2(n397), .C1(n374), 
        .C2(n393), .ZN(n2600) );
  XOR2_X2 U1702 ( .A(n2567), .B(n271), .Z(n1986) );
  OAI21_X4 U1703 ( .B1(n2839), .B2(n345), .A(n2601), .ZN(n2567) );
  AOI222_X2 U1704 ( .A1(n297), .A2(n397), .B1(n319), .B2(n393), .C1(n374), 
        .C2(n390), .ZN(n2601) );
  XOR2_X2 U1705 ( .A(n2568), .B(n271), .Z(n1987) );
  OAI21_X4 U1706 ( .B1(n2840), .B2(n345), .A(n2602), .ZN(n2568) );
  AND2_X4 U1711 ( .A1(n297), .A2(n390), .ZN(n1397) );
  XOR2_X2 U1713 ( .A(n2604), .B(n268), .Z(n1990) );
  OAI21_X4 U1714 ( .B1(n2808), .B2(n342), .A(n2638), .ZN(n2604) );
  NAND2_X4 U1715 ( .A1(n372), .A2(n484), .ZN(n2638) );
  XOR2_X2 U1716 ( .A(n2605), .B(n268), .Z(n1991) );
  OAI21_X4 U1717 ( .B1(n2809), .B2(n342), .A(n2639), .ZN(n2605) );
  AOI21_X4 U1718 ( .B1(n372), .B2(n481), .A(n1398), .ZN(n2639) );
  AND2_X4 U1719 ( .A1(n317), .A2(n484), .ZN(n1398) );
  XOR2_X2 U1720 ( .A(n2606), .B(n268), .Z(n1992) );
  OAI21_X4 U1721 ( .B1(n2810), .B2(n342), .A(n2640), .ZN(n2606) );
  AOI222_X2 U1722 ( .A1(n295), .A2(n484), .B1(n317), .B2(n481), .C1(n372), 
        .C2(n478), .ZN(n2640) );
  XOR2_X2 U1723 ( .A(n2607), .B(n268), .Z(n1993) );
  OAI21_X4 U1724 ( .B1(n2811), .B2(n342), .A(n2641), .ZN(n2607) );
  AOI222_X2 U1725 ( .A1(n295), .A2(n481), .B1(n317), .B2(n478), .C1(n372), 
        .C2(n475), .ZN(n2641) );
  XOR2_X2 U1726 ( .A(n2608), .B(n268), .Z(n1994) );
  OAI21_X4 U1727 ( .B1(n2812), .B2(n342), .A(n2642), .ZN(n2608) );
  AOI222_X2 U1728 ( .A1(n295), .A2(n478), .B1(n317), .B2(n475), .C1(n372), 
        .C2(n472), .ZN(n2642) );
  XOR2_X2 U1729 ( .A(n2609), .B(n268), .Z(n1995) );
  OAI21_X4 U1730 ( .B1(n2813), .B2(n342), .A(n2643), .ZN(n2609) );
  AOI222_X2 U1731 ( .A1(n295), .A2(n475), .B1(n317), .B2(n472), .C1(n372), 
        .C2(n469), .ZN(n2643) );
  XOR2_X2 U1732 ( .A(n2610), .B(n268), .Z(n1996) );
  OAI21_X4 U1733 ( .B1(n2814), .B2(n342), .A(n2644), .ZN(n2610) );
  AOI222_X2 U1734 ( .A1(n295), .A2(n472), .B1(n317), .B2(n469), .C1(n372), 
        .C2(n466), .ZN(n2644) );
  XOR2_X2 U1735 ( .A(n2611), .B(n268), .Z(n1997) );
  OAI21_X4 U1736 ( .B1(n2815), .B2(n342), .A(n2645), .ZN(n2611) );
  AOI222_X2 U1737 ( .A1(n295), .A2(n469), .B1(n317), .B2(n466), .C1(n372), 
        .C2(n463), .ZN(n2645) );
  XOR2_X2 U1738 ( .A(n2612), .B(n268), .Z(n1998) );
  OAI21_X4 U1739 ( .B1(n2816), .B2(n342), .A(n2646), .ZN(n2612) );
  AOI222_X2 U1740 ( .A1(n295), .A2(n466), .B1(n317), .B2(n463), .C1(n372), 
        .C2(n460), .ZN(n2646) );
  XOR2_X2 U1741 ( .A(n2613), .B(n268), .Z(n1999) );
  OAI21_X4 U1742 ( .B1(n2817), .B2(n342), .A(n2647), .ZN(n2613) );
  AOI222_X2 U1743 ( .A1(n295), .A2(n463), .B1(n317), .B2(n460), .C1(n372), 
        .C2(n457), .ZN(n2647) );
  XOR2_X2 U1744 ( .A(n2614), .B(n268), .Z(n2000) );
  OAI21_X4 U1745 ( .B1(n2818), .B2(n342), .A(n2648), .ZN(n2614) );
  AOI222_X2 U1746 ( .A1(n295), .A2(n460), .B1(n317), .B2(n457), .C1(n372), 
        .C2(n454), .ZN(n2648) );
  XOR2_X2 U1747 ( .A(n2615), .B(n268), .Z(n2001) );
  OAI21_X4 U1748 ( .B1(n2819), .B2(n342), .A(n2649), .ZN(n2615) );
  AOI222_X2 U1749 ( .A1(n295), .A2(n457), .B1(n317), .B2(n454), .C1(n372), 
        .C2(n451), .ZN(n2649) );
  XOR2_X2 U1750 ( .A(n2616), .B(n268), .Z(n2002) );
  OAI21_X4 U1751 ( .B1(n2820), .B2(n342), .A(n2650), .ZN(n2616) );
  AOI222_X2 U1752 ( .A1(n295), .A2(n454), .B1(n317), .B2(n451), .C1(n372), 
        .C2(n448), .ZN(n2650) );
  XOR2_X2 U1753 ( .A(n2617), .B(n268), .Z(n2003) );
  OAI21_X4 U1754 ( .B1(n2821), .B2(n342), .A(n2651), .ZN(n2617) );
  AOI222_X2 U1755 ( .A1(n295), .A2(n451), .B1(n317), .B2(n448), .C1(n372), 
        .C2(n445), .ZN(n2651) );
  XOR2_X2 U1756 ( .A(n2618), .B(n268), .Z(n2004) );
  OAI21_X4 U1757 ( .B1(n2822), .B2(n342), .A(n2652), .ZN(n2618) );
  AOI222_X2 U1758 ( .A1(n295), .A2(n448), .B1(n317), .B2(n445), .C1(n372), 
        .C2(n442), .ZN(n2652) );
  XOR2_X2 U1759 ( .A(n2619), .B(n268), .Z(n2005) );
  OAI21_X4 U1760 ( .B1(n2823), .B2(n342), .A(n2653), .ZN(n2619) );
  AOI222_X2 U1761 ( .A1(n295), .A2(n445), .B1(n317), .B2(n442), .C1(n372), 
        .C2(n439), .ZN(n2653) );
  XOR2_X2 U1762 ( .A(n2620), .B(n268), .Z(n2006) );
  OAI21_X4 U1763 ( .B1(n2824), .B2(n342), .A(n2654), .ZN(n2620) );
  AOI222_X2 U1764 ( .A1(n295), .A2(n442), .B1(n317), .B2(n439), .C1(n372), 
        .C2(n436), .ZN(n2654) );
  XOR2_X2 U1765 ( .A(n2621), .B(n268), .Z(n2007) );
  OAI21_X4 U1766 ( .B1(n2825), .B2(n342), .A(n2655), .ZN(n2621) );
  AOI222_X2 U1767 ( .A1(n295), .A2(n439), .B1(n317), .B2(n436), .C1(n372), 
        .C2(n433), .ZN(n2655) );
  XOR2_X2 U1768 ( .A(n2622), .B(n268), .Z(n2008) );
  OAI21_X4 U1769 ( .B1(n2826), .B2(n342), .A(n2656), .ZN(n2622) );
  AOI222_X2 U1770 ( .A1(n295), .A2(n436), .B1(n317), .B2(n433), .C1(n372), 
        .C2(n430), .ZN(n2656) );
  XOR2_X2 U1771 ( .A(n2623), .B(n268), .Z(n2009) );
  OAI21_X4 U1772 ( .B1(n2827), .B2(n342), .A(n2657), .ZN(n2623) );
  AOI222_X2 U1773 ( .A1(n295), .A2(n433), .B1(n317), .B2(n430), .C1(n372), 
        .C2(n427), .ZN(n2657) );
  XOR2_X2 U1774 ( .A(n2624), .B(n268), .Z(n2010) );
  OAI21_X4 U1775 ( .B1(n2828), .B2(n342), .A(n2658), .ZN(n2624) );
  AOI222_X2 U1776 ( .A1(n295), .A2(n430), .B1(n317), .B2(n427), .C1(n372), 
        .C2(n424), .ZN(n2658) );
  XOR2_X2 U1777 ( .A(n2625), .B(n268), .Z(n2011) );
  OAI21_X4 U1778 ( .B1(n2829), .B2(n342), .A(n2659), .ZN(n2625) );
  AOI222_X2 U1779 ( .A1(n295), .A2(n427), .B1(n317), .B2(n424), .C1(n372), 
        .C2(n421), .ZN(n2659) );
  XOR2_X2 U1780 ( .A(n2626), .B(n268), .Z(n2012) );
  OAI21_X4 U1781 ( .B1(n2830), .B2(n342), .A(n2660), .ZN(n2626) );
  AOI222_X2 U1782 ( .A1(n295), .A2(n424), .B1(n317), .B2(n421), .C1(n372), 
        .C2(n418), .ZN(n2660) );
  XOR2_X2 U1783 ( .A(n2627), .B(n268), .Z(n2013) );
  OAI21_X4 U1784 ( .B1(n2831), .B2(n342), .A(n2661), .ZN(n2627) );
  AOI222_X2 U1785 ( .A1(n295), .A2(n421), .B1(n317), .B2(n418), .C1(n372), 
        .C2(n415), .ZN(n2661) );
  XOR2_X2 U1786 ( .A(n2628), .B(n268), .Z(n2014) );
  OAI21_X4 U1787 ( .B1(n2832), .B2(n342), .A(n2662), .ZN(n2628) );
  AOI222_X2 U1788 ( .A1(n295), .A2(n418), .B1(n317), .B2(n415), .C1(n372), 
        .C2(n412), .ZN(n2662) );
  XOR2_X2 U1789 ( .A(n2629), .B(n268), .Z(n2015) );
  OAI21_X4 U1790 ( .B1(n2833), .B2(n342), .A(n2663), .ZN(n2629) );
  AOI222_X2 U1791 ( .A1(n295), .A2(n415), .B1(n317), .B2(n412), .C1(n372), 
        .C2(n409), .ZN(n2663) );
  XOR2_X2 U1792 ( .A(n2630), .B(n268), .Z(n2016) );
  OAI21_X4 U1793 ( .B1(n2834), .B2(n342), .A(n2664), .ZN(n2630) );
  AOI222_X2 U1794 ( .A1(n295), .A2(n412), .B1(n317), .B2(n409), .C1(n372), 
        .C2(n406), .ZN(n2664) );
  XOR2_X2 U1795 ( .A(n2631), .B(n268), .Z(n2017) );
  OAI21_X4 U1796 ( .B1(n2835), .B2(n342), .A(n2665), .ZN(n2631) );
  AOI222_X2 U1797 ( .A1(n295), .A2(n409), .B1(n317), .B2(n406), .C1(n372), 
        .C2(n403), .ZN(n2665) );
  XOR2_X2 U1798 ( .A(n2632), .B(n268), .Z(n2018) );
  OAI21_X4 U1799 ( .B1(n2836), .B2(n342), .A(n2666), .ZN(n2632) );
  AOI222_X2 U1800 ( .A1(n295), .A2(n406), .B1(n317), .B2(n403), .C1(n372), 
        .C2(n400), .ZN(n2666) );
  XOR2_X2 U1801 ( .A(n2633), .B(n268), .Z(n2019) );
  OAI21_X4 U1802 ( .B1(n2837), .B2(n342), .A(n2667), .ZN(n2633) );
  AOI222_X2 U1803 ( .A1(n295), .A2(n403), .B1(n317), .B2(n400), .C1(n372), 
        .C2(n397), .ZN(n2667) );
  XOR2_X2 U1804 ( .A(n2634), .B(n268), .Z(n2020) );
  OAI21_X4 U1805 ( .B1(n2838), .B2(n342), .A(n2668), .ZN(n2634) );
  AOI222_X2 U1806 ( .A1(n295), .A2(n400), .B1(n317), .B2(n397), .C1(n372), 
        .C2(n393), .ZN(n2668) );
  XOR2_X2 U1807 ( .A(n2635), .B(n268), .Z(n2021) );
  AND2_X4 U1816 ( .A1(n295), .A2(n390), .ZN(n1400) );
  XOR2_X2 U1818 ( .A(n2672), .B(n265), .Z(n2025) );
  OAI21_X4 U1819 ( .B1(n2808), .B2(n3127), .A(n2706), .ZN(n2672) );
  NAND2_X4 U1820 ( .A1(n370), .A2(n484), .ZN(n2706) );
  XOR2_X2 U1821 ( .A(n2673), .B(n265), .Z(n2026) );
  OAI21_X4 U1822 ( .B1(n2809), .B2(n339), .A(n2707), .ZN(n2673) );
  AOI21_X4 U1823 ( .B1(n370), .B2(n481), .A(n1401), .ZN(n2707) );
  AND2_X4 U1824 ( .A1(n315), .A2(n484), .ZN(n1401) );
  XOR2_X2 U1825 ( .A(n2674), .B(n265), .Z(n2027) );
  OAI21_X4 U1826 ( .B1(n2810), .B2(n3127), .A(n2708), .ZN(n2674) );
  AOI222_X2 U1827 ( .A1(n293), .A2(n484), .B1(n315), .B2(n481), .C1(n370), 
        .C2(n478), .ZN(n2708) );
  XOR2_X2 U1828 ( .A(n2675), .B(n265), .Z(n2028) );
  OAI21_X4 U1829 ( .B1(n2811), .B2(n339), .A(n2709), .ZN(n2675) );
  AOI222_X2 U1830 ( .A1(n293), .A2(n481), .B1(n315), .B2(n478), .C1(n370), 
        .C2(n475), .ZN(n2709) );
  XOR2_X2 U1831 ( .A(n2676), .B(n265), .Z(n2029) );
  OAI21_X4 U1832 ( .B1(n2812), .B2(n339), .A(n2710), .ZN(n2676) );
  AOI222_X2 U1833 ( .A1(n293), .A2(n478), .B1(n315), .B2(n475), .C1(n370), 
        .C2(n472), .ZN(n2710) );
  XOR2_X2 U1834 ( .A(n2677), .B(n265), .Z(n2030) );
  OAI21_X4 U1835 ( .B1(n2813), .B2(n339), .A(n2711), .ZN(n2677) );
  AOI222_X2 U1836 ( .A1(n293), .A2(n475), .B1(n315), .B2(n472), .C1(n370), 
        .C2(n469), .ZN(n2711) );
  XOR2_X2 U1837 ( .A(n2678), .B(n265), .Z(n2031) );
  OAI21_X4 U1838 ( .B1(n2814), .B2(n339), .A(n2712), .ZN(n2678) );
  AOI222_X2 U1839 ( .A1(n293), .A2(n472), .B1(n315), .B2(n469), .C1(n370), 
        .C2(n466), .ZN(n2712) );
  XOR2_X2 U1840 ( .A(n2679), .B(n265), .Z(n2032) );
  OAI21_X4 U1841 ( .B1(n2815), .B2(n339), .A(n2713), .ZN(n2679) );
  AOI222_X2 U1842 ( .A1(n293), .A2(n469), .B1(n315), .B2(n466), .C1(n370), 
        .C2(n463), .ZN(n2713) );
  XOR2_X2 U1843 ( .A(n2680), .B(n265), .Z(n2033) );
  OAI21_X4 U1844 ( .B1(n2816), .B2(n339), .A(n2714), .ZN(n2680) );
  AOI222_X2 U1845 ( .A1(n293), .A2(n466), .B1(n315), .B2(n463), .C1(n370), 
        .C2(n460), .ZN(n2714) );
  XOR2_X2 U1846 ( .A(n2681), .B(n265), .Z(n2034) );
  OAI21_X4 U1847 ( .B1(n2817), .B2(n339), .A(n2715), .ZN(n2681) );
  AOI222_X2 U1848 ( .A1(n293), .A2(n463), .B1(n315), .B2(n460), .C1(n370), 
        .C2(n457), .ZN(n2715) );
  XOR2_X2 U1849 ( .A(n2682), .B(n265), .Z(n2035) );
  OAI21_X4 U1850 ( .B1(n2818), .B2(n339), .A(n2716), .ZN(n2682) );
  AOI222_X2 U1851 ( .A1(n293), .A2(n460), .B1(n315), .B2(n457), .C1(n370), 
        .C2(n454), .ZN(n2716) );
  XOR2_X2 U1852 ( .A(n2683), .B(n265), .Z(n2036) );
  OAI21_X4 U1853 ( .B1(n2819), .B2(n339), .A(n2717), .ZN(n2683) );
  AOI222_X2 U1854 ( .A1(n293), .A2(n457), .B1(n315), .B2(n454), .C1(n370), 
        .C2(n451), .ZN(n2717) );
  XOR2_X2 U1855 ( .A(n2684), .B(n265), .Z(n2037) );
  OAI21_X4 U1856 ( .B1(n2820), .B2(n339), .A(n2718), .ZN(n2684) );
  AOI222_X2 U1857 ( .A1(n293), .A2(n454), .B1(n315), .B2(n451), .C1(n370), 
        .C2(n448), .ZN(n2718) );
  XOR2_X2 U1858 ( .A(n2685), .B(n265), .Z(n2038) );
  OAI21_X4 U1859 ( .B1(n2821), .B2(n339), .A(n2719), .ZN(n2685) );
  AOI222_X2 U1860 ( .A1(n293), .A2(n451), .B1(n315), .B2(n448), .C1(n370), 
        .C2(n445), .ZN(n2719) );
  XOR2_X2 U1861 ( .A(n2686), .B(n265), .Z(n2039) );
  OAI21_X4 U1862 ( .B1(n2822), .B2(n339), .A(n2720), .ZN(n2686) );
  AOI222_X2 U1863 ( .A1(n293), .A2(n448), .B1(n315), .B2(n445), .C1(n370), 
        .C2(n442), .ZN(n2720) );
  XOR2_X2 U1864 ( .A(n2687), .B(n265), .Z(n2040) );
  OAI21_X4 U1865 ( .B1(n2823), .B2(n339), .A(n2721), .ZN(n2687) );
  AOI222_X2 U1866 ( .A1(n293), .A2(n445), .B1(n315), .B2(n442), .C1(n370), 
        .C2(n439), .ZN(n2721) );
  XOR2_X2 U1867 ( .A(n2688), .B(n265), .Z(n2041) );
  OAI21_X4 U1868 ( .B1(n2824), .B2(n339), .A(n2722), .ZN(n2688) );
  AOI222_X2 U1869 ( .A1(n293), .A2(n442), .B1(n315), .B2(n439), .C1(n370), 
        .C2(n436), .ZN(n2722) );
  XOR2_X2 U1870 ( .A(n2689), .B(n265), .Z(n2042) );
  OAI21_X4 U1871 ( .B1(n2825), .B2(n339), .A(n2723), .ZN(n2689) );
  AOI222_X2 U1872 ( .A1(n293), .A2(n439), .B1(n315), .B2(n436), .C1(n370), 
        .C2(n433), .ZN(n2723) );
  XOR2_X2 U1873 ( .A(n2690), .B(n265), .Z(n2043) );
  OAI21_X4 U1874 ( .B1(n2826), .B2(n339), .A(n2724), .ZN(n2690) );
  AOI222_X2 U1875 ( .A1(n293), .A2(n436), .B1(n315), .B2(n433), .C1(n370), 
        .C2(n430), .ZN(n2724) );
  XOR2_X2 U1876 ( .A(n2691), .B(n265), .Z(n2044) );
  OAI21_X4 U1877 ( .B1(n2827), .B2(n339), .A(n2725), .ZN(n2691) );
  AOI222_X2 U1878 ( .A1(n293), .A2(n433), .B1(n315), .B2(n430), .C1(n370), 
        .C2(n427), .ZN(n2725) );
  XOR2_X2 U1879 ( .A(n2692), .B(n265), .Z(n2045) );
  OAI21_X4 U1880 ( .B1(n2828), .B2(n339), .A(n2726), .ZN(n2692) );
  AOI222_X2 U1881 ( .A1(n293), .A2(n430), .B1(n315), .B2(n427), .C1(n370), 
        .C2(n424), .ZN(n2726) );
  XOR2_X2 U1882 ( .A(n2693), .B(n265), .Z(n2046) );
  OAI21_X4 U1883 ( .B1(n2829), .B2(n339), .A(n2727), .ZN(n2693) );
  AOI222_X2 U1884 ( .A1(n293), .A2(n427), .B1(n315), .B2(n424), .C1(n370), 
        .C2(n421), .ZN(n2727) );
  XOR2_X2 U1885 ( .A(n2694), .B(n265), .Z(n2047) );
  OAI21_X4 U1886 ( .B1(n2830), .B2(n339), .A(n2728), .ZN(n2694) );
  AOI222_X2 U1887 ( .A1(n293), .A2(n424), .B1(n315), .B2(n421), .C1(n370), 
        .C2(n418), .ZN(n2728) );
  XOR2_X2 U1888 ( .A(n2695), .B(n265), .Z(n2048) );
  OAI21_X4 U1889 ( .B1(n2831), .B2(n339), .A(n2729), .ZN(n2695) );
  AOI222_X2 U1890 ( .A1(n293), .A2(n421), .B1(n315), .B2(n418), .C1(n370), 
        .C2(n415), .ZN(n2729) );
  XOR2_X2 U1891 ( .A(n2696), .B(n265), .Z(n2049) );
  OAI21_X4 U1892 ( .B1(n2832), .B2(n339), .A(n2730), .ZN(n2696) );
  AOI222_X2 U1893 ( .A1(n293), .A2(n418), .B1(n315), .B2(n415), .C1(n370), 
        .C2(n412), .ZN(n2730) );
  XOR2_X2 U1894 ( .A(n2697), .B(n265), .Z(n2050) );
  OAI21_X4 U1895 ( .B1(n2833), .B2(n339), .A(n2731), .ZN(n2697) );
  AOI222_X2 U1896 ( .A1(n293), .A2(n415), .B1(n315), .B2(n412), .C1(n370), 
        .C2(n409), .ZN(n2731) );
  XOR2_X2 U1897 ( .A(n2698), .B(n265), .Z(n2051) );
  OAI21_X4 U1898 ( .B1(n2834), .B2(n339), .A(n2732), .ZN(n2698) );
  AOI222_X2 U1899 ( .A1(n293), .A2(n412), .B1(n315), .B2(n409), .C1(n370), 
        .C2(n406), .ZN(n2732) );
  XOR2_X2 U1900 ( .A(n2699), .B(n265), .Z(n2052) );
  OAI21_X4 U1901 ( .B1(n2835), .B2(n339), .A(n2733), .ZN(n2699) );
  AOI222_X2 U1902 ( .A1(n293), .A2(n409), .B1(n315), .B2(n406), .C1(n370), 
        .C2(n403), .ZN(n2733) );
  XOR2_X2 U1903 ( .A(n2700), .B(n265), .Z(n2053) );
  OAI21_X4 U1904 ( .B1(n2836), .B2(n339), .A(n2734), .ZN(n2700) );
  AOI222_X2 U1905 ( .A1(n293), .A2(n406), .B1(n315), .B2(n403), .C1(n370), 
        .C2(n400), .ZN(n2734) );
  XOR2_X2 U1906 ( .A(n2701), .B(n265), .Z(n2054) );
  OAI21_X4 U1907 ( .B1(n2837), .B2(n339), .A(n2735), .ZN(n2701) );
  AOI222_X2 U1908 ( .A1(n293), .A2(n403), .B1(n315), .B2(n400), .C1(n370), 
        .C2(n397), .ZN(n2735) );
  XOR2_X2 U1909 ( .A(n2702), .B(n265), .Z(n2055) );
  OAI21_X4 U1910 ( .B1(n2838), .B2(n339), .A(n2736), .ZN(n2702) );
  AOI222_X2 U1911 ( .A1(n293), .A2(n400), .B1(n315), .B2(n397), .C1(n370), 
        .C2(n393), .ZN(n2736) );
  XOR2_X2 U1912 ( .A(n2703), .B(n265), .Z(n2056) );
  OAI21_X4 U1913 ( .B1(n2839), .B2(n339), .A(n2737), .ZN(n2703) );
  AOI222_X2 U1914 ( .A1(n293), .A2(n397), .B1(n315), .B2(n393), .C1(n370), 
        .C2(n390), .ZN(n2737) );
  XOR2_X2 U1915 ( .A(n2704), .B(n265), .Z(n2057) );
  OAI21_X4 U1916 ( .B1(n2840), .B2(n339), .A(n2738), .ZN(n2704) );
  OAI21_X4 U1919 ( .B1(n2841), .B2(n339), .A(n2739), .ZN(n2705) );
  AND2_X4 U1921 ( .A1(n293), .A2(n390), .ZN(n1403) );
  XOR2_X2 U1923 ( .A(n2740), .B(n262), .Z(n2060) );
  OAI21_X4 U1924 ( .B1(n2808), .B2(n3126), .A(n2774), .ZN(n2740) );
  NAND2_X4 U1925 ( .A1(n368), .A2(n484), .ZN(n2774) );
  XOR2_X2 U1926 ( .A(n2741), .B(n262), .Z(n2061) );
  OAI21_X4 U1927 ( .B1(n2809), .B2(n3126), .A(n2775), .ZN(n2741) );
  AOI21_X4 U1928 ( .B1(n368), .B2(n481), .A(n1404), .ZN(n2775) );
  AND2_X4 U1929 ( .A1(n313), .A2(n484), .ZN(n1404) );
  XOR2_X2 U1930 ( .A(n2742), .B(n262), .Z(n2062) );
  OAI21_X4 U1931 ( .B1(n2810), .B2(n3126), .A(n2776), .ZN(n2742) );
  AOI222_X2 U1932 ( .A1(n3226), .A2(n484), .B1(n313), .B2(n481), .C1(n368), 
        .C2(n478), .ZN(n2776) );
  XOR2_X2 U1933 ( .A(n2743), .B(n262), .Z(n2063) );
  OAI21_X4 U1934 ( .B1(n2811), .B2(n336), .A(n2777), .ZN(n2743) );
  AOI222_X2 U1935 ( .A1(n3226), .A2(n481), .B1(n313), .B2(n478), .C1(n368), 
        .C2(n475), .ZN(n2777) );
  XOR2_X2 U1936 ( .A(n2744), .B(n262), .Z(n2064) );
  OAI21_X4 U1937 ( .B1(n2812), .B2(n336), .A(n2778), .ZN(n2744) );
  AOI222_X2 U1938 ( .A1(n3226), .A2(n478), .B1(n313), .B2(n475), .C1(n368), 
        .C2(n472), .ZN(n2778) );
  XOR2_X2 U1939 ( .A(n2745), .B(n262), .Z(n2065) );
  OAI21_X4 U1940 ( .B1(n2813), .B2(n336), .A(n2779), .ZN(n2745) );
  AOI222_X2 U1941 ( .A1(n3226), .A2(n475), .B1(n313), .B2(n472), .C1(n368), 
        .C2(n469), .ZN(n2779) );
  XOR2_X2 U1942 ( .A(n2746), .B(n262), .Z(n2066) );
  OAI21_X4 U1943 ( .B1(n2814), .B2(n336), .A(n2780), .ZN(n2746) );
  AOI222_X2 U1944 ( .A1(n3226), .A2(n472), .B1(n313), .B2(n469), .C1(n368), 
        .C2(n466), .ZN(n2780) );
  XOR2_X2 U1945 ( .A(n2747), .B(n262), .Z(n2067) );
  OAI21_X4 U1946 ( .B1(n2815), .B2(n336), .A(n2781), .ZN(n2747) );
  AOI222_X2 U1947 ( .A1(n3226), .A2(n469), .B1(n313), .B2(n466), .C1(n368), 
        .C2(n463), .ZN(n2781) );
  XOR2_X2 U1948 ( .A(n2748), .B(n262), .Z(n2068) );
  OAI21_X4 U1949 ( .B1(n2816), .B2(n336), .A(n2782), .ZN(n2748) );
  AOI222_X2 U1950 ( .A1(n3226), .A2(n466), .B1(n313), .B2(n463), .C1(n368), 
        .C2(n460), .ZN(n2782) );
  XOR2_X2 U1951 ( .A(n2749), .B(n262), .Z(n2069) );
  OAI21_X4 U1952 ( .B1(n2817), .B2(n336), .A(n2783), .ZN(n2749) );
  AOI222_X2 U1953 ( .A1(n3226), .A2(n463), .B1(n313), .B2(n460), .C1(n368), 
        .C2(n457), .ZN(n2783) );
  XOR2_X2 U1954 ( .A(n2750), .B(n262), .Z(n2070) );
  OAI21_X4 U1955 ( .B1(n2818), .B2(n336), .A(n2784), .ZN(n2750) );
  AOI222_X2 U1956 ( .A1(n3226), .A2(n460), .B1(n313), .B2(n457), .C1(n368), 
        .C2(n454), .ZN(n2784) );
  XOR2_X2 U1957 ( .A(n2751), .B(n262), .Z(n2071) );
  OAI21_X4 U1958 ( .B1(n2819), .B2(n336), .A(n2785), .ZN(n2751) );
  AOI222_X2 U1959 ( .A1(n3226), .A2(n457), .B1(n313), .B2(n454), .C1(n368), 
        .C2(n451), .ZN(n2785) );
  XOR2_X2 U1960 ( .A(n2752), .B(n262), .Z(n2072) );
  OAI21_X4 U1961 ( .B1(n2820), .B2(n336), .A(n2786), .ZN(n2752) );
  AOI222_X2 U1962 ( .A1(n3226), .A2(n454), .B1(n313), .B2(n451), .C1(n368), 
        .C2(n448), .ZN(n2786) );
  XOR2_X2 U1963 ( .A(n2753), .B(n262), .Z(n2073) );
  OAI21_X4 U1964 ( .B1(n2821), .B2(n336), .A(n2787), .ZN(n2753) );
  AOI222_X2 U1965 ( .A1(n3226), .A2(n451), .B1(n313), .B2(n448), .C1(n368), 
        .C2(n445), .ZN(n2787) );
  XOR2_X2 U1966 ( .A(n2754), .B(n262), .Z(n2074) );
  OAI21_X4 U1967 ( .B1(n2822), .B2(n336), .A(n2788), .ZN(n2754) );
  AOI222_X2 U1968 ( .A1(n3226), .A2(n448), .B1(n313), .B2(n445), .C1(n368), 
        .C2(n442), .ZN(n2788) );
  XOR2_X2 U1969 ( .A(n2755), .B(n262), .Z(n2075) );
  OAI21_X4 U1970 ( .B1(n2823), .B2(n336), .A(n2789), .ZN(n2755) );
  AOI222_X2 U1971 ( .A1(n3226), .A2(n445), .B1(n313), .B2(n442), .C1(n368), 
        .C2(n439), .ZN(n2789) );
  XOR2_X2 U1972 ( .A(n2756), .B(n262), .Z(n2076) );
  OAI21_X4 U1973 ( .B1(n2824), .B2(n336), .A(n2790), .ZN(n2756) );
  AOI222_X2 U1974 ( .A1(n3226), .A2(n442), .B1(n313), .B2(n439), .C1(n368), 
        .C2(n436), .ZN(n2790) );
  XOR2_X2 U1975 ( .A(n2757), .B(n262), .Z(n2077) );
  OAI21_X4 U1976 ( .B1(n2825), .B2(n336), .A(n2791), .ZN(n2757) );
  AOI222_X2 U1977 ( .A1(n3226), .A2(n439), .B1(n313), .B2(n436), .C1(n368), 
        .C2(n433), .ZN(n2791) );
  XOR2_X2 U1978 ( .A(n2758), .B(n262), .Z(n2078) );
  OAI21_X4 U1979 ( .B1(n2826), .B2(n336), .A(n2792), .ZN(n2758) );
  AOI222_X2 U1980 ( .A1(n3226), .A2(n436), .B1(n313), .B2(n433), .C1(n368), 
        .C2(n430), .ZN(n2792) );
  XOR2_X2 U1981 ( .A(n2759), .B(n262), .Z(n2079) );
  OAI21_X4 U1982 ( .B1(n2827), .B2(n336), .A(n2793), .ZN(n2759) );
  AOI222_X2 U1983 ( .A1(n3226), .A2(n433), .B1(n313), .B2(n430), .C1(n368), 
        .C2(n427), .ZN(n2793) );
  XOR2_X2 U1984 ( .A(n2760), .B(n262), .Z(n2080) );
  OAI21_X4 U1985 ( .B1(n2828), .B2(n336), .A(n2794), .ZN(n2760) );
  AOI222_X2 U1986 ( .A1(n3226), .A2(n430), .B1(n313), .B2(n427), .C1(n368), 
        .C2(n424), .ZN(n2794) );
  XOR2_X2 U1987 ( .A(n2761), .B(n262), .Z(n2081) );
  OAI21_X4 U1988 ( .B1(n2829), .B2(n336), .A(n2795), .ZN(n2761) );
  AOI222_X2 U1989 ( .A1(n3226), .A2(n427), .B1(n313), .B2(n424), .C1(n368), 
        .C2(n421), .ZN(n2795) );
  XOR2_X2 U1990 ( .A(n2762), .B(n262), .Z(n2082) );
  OAI21_X4 U1991 ( .B1(n2830), .B2(n336), .A(n2796), .ZN(n2762) );
  AOI222_X2 U1992 ( .A1(n3226), .A2(n424), .B1(n313), .B2(n421), .C1(n368), 
        .C2(n418), .ZN(n2796) );
  XOR2_X2 U1993 ( .A(n2763), .B(n262), .Z(n2083) );
  OAI21_X4 U1994 ( .B1(n2831), .B2(n336), .A(n2797), .ZN(n2763) );
  AOI222_X2 U1995 ( .A1(n3226), .A2(n421), .B1(n313), .B2(n418), .C1(n368), 
        .C2(n415), .ZN(n2797) );
  XOR2_X2 U1996 ( .A(n2764), .B(n262), .Z(n2084) );
  OAI21_X4 U1997 ( .B1(n2832), .B2(n336), .A(n2798), .ZN(n2764) );
  AOI222_X2 U1998 ( .A1(n3226), .A2(n418), .B1(n313), .B2(n415), .C1(n368), 
        .C2(n412), .ZN(n2798) );
  XOR2_X2 U1999 ( .A(n2765), .B(n262), .Z(n2085) );
  OAI21_X4 U2000 ( .B1(n2833), .B2(n336), .A(n2799), .ZN(n2765) );
  AOI222_X2 U2001 ( .A1(n3226), .A2(n415), .B1(n313), .B2(n412), .C1(n368), 
        .C2(n409), .ZN(n2799) );
  XOR2_X2 U2002 ( .A(n2766), .B(n262), .Z(n2086) );
  OAI21_X4 U2003 ( .B1(n2834), .B2(n336), .A(n2800), .ZN(n2766) );
  AOI222_X2 U2004 ( .A1(n3226), .A2(n412), .B1(n313), .B2(n409), .C1(n368), 
        .C2(n406), .ZN(n2800) );
  XOR2_X2 U2005 ( .A(n2767), .B(n262), .Z(n2087) );
  OAI21_X4 U2006 ( .B1(n2835), .B2(n336), .A(n2801), .ZN(n2767) );
  AOI222_X2 U2007 ( .A1(n3226), .A2(n409), .B1(n313), .B2(n406), .C1(n368), 
        .C2(n403), .ZN(n2801) );
  XOR2_X2 U2008 ( .A(n2768), .B(n262), .Z(n2088) );
  OAI21_X4 U2009 ( .B1(n2836), .B2(n336), .A(n2802), .ZN(n2768) );
  AOI222_X2 U2010 ( .A1(n3226), .A2(n406), .B1(n313), .B2(n403), .C1(n368), 
        .C2(n400), .ZN(n2802) );
  XOR2_X2 U2011 ( .A(n2769), .B(n262), .Z(n2089) );
  OAI21_X4 U2012 ( .B1(n2837), .B2(n336), .A(n2803), .ZN(n2769) );
  AOI222_X2 U2013 ( .A1(n3226), .A2(n403), .B1(n313), .B2(n400), .C1(n368), 
        .C2(n397), .ZN(n2803) );
  XOR2_X2 U2014 ( .A(n2770), .B(n262), .Z(n2090) );
  OAI21_X4 U2015 ( .B1(n2838), .B2(n336), .A(n2804), .ZN(n2770) );
  AOI222_X2 U2016 ( .A1(n3226), .A2(n400), .B1(n313), .B2(n397), .C1(n368), 
        .C2(n393), .ZN(n2804) );
  XOR2_X2 U2017 ( .A(n2771), .B(n262), .Z(n2091) );
  OAI21_X4 U2018 ( .B1(n2839), .B2(n336), .A(n2805), .ZN(n2771) );
  AOI222_X2 U2019 ( .A1(n3226), .A2(n397), .B1(n313), .B2(n393), .C1(n368), 
        .C2(n390), .ZN(n2805) );
  XOR2_X2 U2020 ( .A(n2772), .B(n262), .Z(n678) );
  OAI21_X4 U2021 ( .B1(n2840), .B2(n336), .A(n2806), .ZN(n2772) );
  XOR2_X2 U2023 ( .A(n2773), .B(n262), .Z(n2093) );
  OAI21_X4 U2024 ( .B1(n2841), .B2(n336), .A(n2807), .ZN(n2773) );
  AND2_X4 U2026 ( .A1(n3226), .A2(n390), .ZN(n1406) );
  AND3_X4 U2103 ( .A1(n2908), .A2(n2919), .A3(a[31]), .ZN(n388) );
  AND3_X4 U2107 ( .A1(n2931), .A2(n2909), .A3(n2920), .ZN(n386) );
  AND3_X4 U2112 ( .A1(n2932), .A2(n2910), .A3(n2921), .ZN(n384) );
  AND3_X4 U2117 ( .A1(n2933), .A2(n2911), .A3(n2922), .ZN(n382) );
  AND3_X4 U2122 ( .A1(n2934), .A2(n2912), .A3(n2923), .ZN(n380) );
  AND3_X4 U2127 ( .A1(n2935), .A2(n2913), .A3(n2924), .ZN(n378) );
  AND3_X4 U2132 ( .A1(n2936), .A2(n2914), .A3(n2925), .ZN(n376) );
  AND3_X4 U2137 ( .A1(n2937), .A2(n2915), .A3(n2926), .ZN(n374) );
  AND3_X4 U2142 ( .A1(n2938), .A2(n2916), .A3(n2927), .ZN(n372) );
  AND3_X4 U2147 ( .A1(n2939), .A2(n2917), .A3(n2928), .ZN(n370) );
  XOR2_X2 U2151 ( .A(a[4]), .B(n265), .Z(n2939) );
  AND3_X4 U2152 ( .A1(n2940), .A2(n2929), .A3(n2918), .ZN(n368) );
  XNOR2_X2 U2158 ( .A(n1441), .B(n1440), .ZN(n2843) );
  NAND2_X4 U2159 ( .A1(n1441), .A2(n484), .ZN(n2808) );
  XOR2_X2 U2162 ( .A(n1452), .B(n1407), .Z(n2844) );
  OAI21_X4 U2163 ( .B1(n1600), .B2(n1442), .A(n1443), .ZN(n1441) );
  NAND2_X4 U2164 ( .A1(n1528), .A2(n1444), .ZN(n1442) );
  AOI21_X4 U2165 ( .B1(n1529), .B2(n1444), .A(n1445), .ZN(n1443) );
  NOR2_X4 U2166 ( .A1(n1488), .A2(n1446), .ZN(n1444) );
  OAI21_X4 U2167 ( .B1(n1489), .B2(n1446), .A(n1447), .ZN(n1445) );
  NAND2_X4 U2168 ( .A1(n1468), .A2(n1448), .ZN(n1446) );
  AOI21_X4 U2169 ( .B1(n1448), .B2(n1469), .A(n1449), .ZN(n1447) );
  NOR2_X4 U2170 ( .A1(n1459), .A2(n1450), .ZN(n1448) );
  OAI21_X4 U2171 ( .B1(n1450), .B2(n1462), .A(n1451), .ZN(n1449) );
  NAND2_X4 U2172 ( .A1(n1689), .A2(n1451), .ZN(n1407) );
  NOR2_X4 U2174 ( .A1(n481), .A2(n484), .ZN(n1450) );
  NAND2_X4 U2175 ( .A1(n481), .A2(n484), .ZN(n1451) );
  XOR2_X2 U2176 ( .A(n1463), .B(n1408), .Z(n2845) );
  AOI21_X4 U2177 ( .B1(n1599), .B2(n1453), .A(n1454), .ZN(n1452) );
  NOR2_X4 U2178 ( .A1(n1530), .A2(n1455), .ZN(n1453) );
  OAI21_X4 U2179 ( .B1(n1531), .B2(n1455), .A(n1456), .ZN(n1454) );
  NAND2_X4 U2180 ( .A1(n1457), .A2(n1490), .ZN(n1455) );
  AOI21_X4 U2181 ( .B1(n1457), .B2(n1491), .A(n1458), .ZN(n1456) );
  NOR2_X4 U2182 ( .A1(n1470), .A2(n1459), .ZN(n1457) );
  OAI21_X4 U2183 ( .B1(n1471), .B2(n1459), .A(n1462), .ZN(n1458) );
  NAND2_X4 U2186 ( .A1(n1690), .A2(n1462), .ZN(n1408) );
  NOR2_X4 U2188 ( .A1(n478), .A2(n481), .ZN(n1459) );
  NAND2_X4 U2189 ( .A1(n478), .A2(n481), .ZN(n1462) );
  XOR2_X2 U2190 ( .A(n1476), .B(n1409), .Z(n2846) );
  AOI21_X4 U2191 ( .B1(n1599), .B2(n1464), .A(n1465), .ZN(n1463) );
  NOR2_X4 U2192 ( .A1(n1530), .A2(n1466), .ZN(n1464) );
  OAI21_X4 U2193 ( .B1(n1531), .B2(n1466), .A(n1467), .ZN(n1465) );
  NAND2_X4 U2194 ( .A1(n1490), .A2(n1468), .ZN(n1466) );
  AOI21_X4 U2195 ( .B1(n1491), .B2(n1468), .A(n1469), .ZN(n1467) );
  NOR2_X4 U2200 ( .A1(n1483), .A2(n1474), .ZN(n1468) );
  OAI21_X4 U2201 ( .B1(n1474), .B2(n1484), .A(n1475), .ZN(n1469) );
  NAND2_X4 U2202 ( .A1(n1691), .A2(n1475), .ZN(n1409) );
  NOR2_X4 U2204 ( .A1(n475), .A2(n478), .ZN(n1474) );
  NAND2_X4 U2205 ( .A1(n475), .A2(n478), .ZN(n1475) );
  XOR2_X2 U2206 ( .A(n1485), .B(n1410), .Z(n2847) );
  AOI21_X4 U2207 ( .B1(n1599), .B2(n1477), .A(n1478), .ZN(n1476) );
  NOR2_X4 U2208 ( .A1(n1530), .A2(n1479), .ZN(n1477) );
  OAI21_X4 U2209 ( .B1(n1531), .B2(n1479), .A(n1480), .ZN(n1478) );
  NAND2_X4 U2210 ( .A1(n1490), .A2(n1692), .ZN(n1479) );
  AOI21_X4 U2211 ( .B1(n1491), .B2(n1692), .A(n1482), .ZN(n1480) );
  NAND2_X4 U2214 ( .A1(n1692), .A2(n1484), .ZN(n1410) );
  NOR2_X4 U2216 ( .A1(n472), .A2(n475), .ZN(n1483) );
  NAND2_X4 U2217 ( .A1(n472), .A2(n475), .ZN(n1484) );
  XOR2_X2 U2218 ( .A(n1498), .B(n1411), .Z(n2848) );
  AOI21_X4 U2219 ( .B1(n1599), .B2(n1486), .A(n1487), .ZN(n1485) );
  NOR2_X4 U2220 ( .A1(n1530), .A2(n1488), .ZN(n1486) );
  OAI21_X4 U2221 ( .B1(n1531), .B2(n1488), .A(n1489), .ZN(n1487) );
  NAND2_X4 U2226 ( .A1(n1512), .A2(n1494), .ZN(n1488) );
  AOI21_X4 U2227 ( .B1(n1494), .B2(n1513), .A(n1495), .ZN(n1489) );
  NOR2_X4 U2228 ( .A1(n1505), .A2(n1496), .ZN(n1494) );
  OAI21_X4 U2229 ( .B1(n1496), .B2(n1506), .A(n1497), .ZN(n1495) );
  NAND2_X4 U2230 ( .A1(n1693), .A2(n1497), .ZN(n1411) );
  NOR2_X4 U2232 ( .A1(n469), .A2(n472), .ZN(n1496) );
  NAND2_X4 U2233 ( .A1(n469), .A2(n472), .ZN(n1497) );
  XOR2_X2 U2234 ( .A(n1507), .B(n1412), .Z(n2849) );
  AOI21_X4 U2235 ( .B1(n1599), .B2(n1499), .A(n1500), .ZN(n1498) );
  NOR2_X4 U2236 ( .A1(n1530), .A2(n1501), .ZN(n1499) );
  OAI21_X4 U2237 ( .B1(n1531), .B2(n1501), .A(n1502), .ZN(n1500) );
  NAND2_X4 U2238 ( .A1(n1512), .A2(n1694), .ZN(n1501) );
  AOI21_X4 U2239 ( .B1(n1513), .B2(n1694), .A(n1504), .ZN(n1502) );
  NAND2_X4 U2242 ( .A1(n1694), .A2(n1506), .ZN(n1412) );
  NOR2_X4 U2244 ( .A1(n466), .A2(n469), .ZN(n1505) );
  NAND2_X4 U2245 ( .A1(n466), .A2(n469), .ZN(n1506) );
  XOR2_X2 U2246 ( .A(n1520), .B(n1413), .Z(n2850) );
  AOI21_X4 U2247 ( .B1(n1599), .B2(n1508), .A(n1509), .ZN(n1507) );
  NOR2_X4 U2248 ( .A1(n1530), .A2(n1510), .ZN(n1508) );
  OAI21_X4 U2249 ( .B1(n1531), .B2(n1510), .A(n1511), .ZN(n1509) );
  NOR2_X4 U2256 ( .A1(n1523), .A2(n1518), .ZN(n1512) );
  OAI21_X4 U2257 ( .B1(n1518), .B2(n1526), .A(n1519), .ZN(n1513) );
  NAND2_X4 U2258 ( .A1(n1695), .A2(n1519), .ZN(n1413) );
  NOR2_X4 U2260 ( .A1(n463), .A2(n466), .ZN(n1518) );
  NAND2_X4 U2261 ( .A1(n463), .A2(n466), .ZN(n1519) );
  XOR2_X2 U2262 ( .A(n1527), .B(n1414), .Z(n2851) );
  AOI21_X4 U2263 ( .B1(n1599), .B2(n1521), .A(n1522), .ZN(n1520) );
  NOR2_X4 U2264 ( .A1(n1530), .A2(n1523), .ZN(n1521) );
  OAI21_X4 U2265 ( .B1(n1531), .B2(n1523), .A(n1526), .ZN(n1522) );
  NAND2_X4 U2268 ( .A1(n1696), .A2(n1526), .ZN(n1414) );
  NOR2_X4 U2270 ( .A1(n460), .A2(n463), .ZN(n1523) );
  NAND2_X4 U2271 ( .A1(n460), .A2(n463), .ZN(n1526) );
  XOR2_X2 U2272 ( .A(n1540), .B(n1415), .Z(n2852) );
  AOI21_X4 U2273 ( .B1(n1599), .B2(n1528), .A(n1529), .ZN(n1527) );
  NOR2_X4 U2278 ( .A1(n1568), .A2(n1534), .ZN(n1528) );
  OAI21_X4 U2279 ( .B1(n1569), .B2(n1534), .A(n1535), .ZN(n1529) );
  NAND2_X4 U2280 ( .A1(n1552), .A2(n1536), .ZN(n1534) );
  AOI21_X4 U2281 ( .B1(n1536), .B2(n1555), .A(n1537), .ZN(n1535) );
  NOR2_X4 U2282 ( .A1(n1543), .A2(n1538), .ZN(n1536) );
  OAI21_X4 U2283 ( .B1(n1538), .B2(n1546), .A(n1539), .ZN(n1537) );
  NAND2_X4 U2284 ( .A1(n1697), .A2(n1539), .ZN(n1415) );
  NOR2_X4 U2286 ( .A1(n457), .A2(n460), .ZN(n1538) );
  NAND2_X4 U2287 ( .A1(n457), .A2(n460), .ZN(n1539) );
  XOR2_X2 U2288 ( .A(n1547), .B(n1416), .Z(n2853) );
  AOI21_X4 U2289 ( .B1(n1599), .B2(n1541), .A(n1542), .ZN(n1540) );
  NOR2_X4 U2290 ( .A1(n1550), .A2(n1543), .ZN(n1541) );
  OAI21_X4 U2291 ( .B1(n1551), .B2(n1543), .A(n1546), .ZN(n1542) );
  NAND2_X4 U2294 ( .A1(n1698), .A2(n1546), .ZN(n1416) );
  NOR2_X4 U2296 ( .A1(n454), .A2(n457), .ZN(n1543) );
  NAND2_X4 U2297 ( .A1(n454), .A2(n457), .ZN(n1546) );
  XOR2_X2 U2298 ( .A(n1558), .B(n1417), .Z(n2854) );
  AOI21_X4 U2299 ( .B1(n1599), .B2(n1548), .A(n1549), .ZN(n1547) );
  NAND2_X4 U2302 ( .A1(n1570), .A2(n1552), .ZN(n1550) );
  AOI21_X4 U2303 ( .B1(n1571), .B2(n1552), .A(n1555), .ZN(n1551) );
  NOR2_X4 U2306 ( .A1(n1561), .A2(n1556), .ZN(n1552) );
  OAI21_X4 U2307 ( .B1(n1556), .B2(n1564), .A(n1557), .ZN(n1555) );
  NAND2_X4 U2308 ( .A1(n1699), .A2(n1557), .ZN(n1417) );
  NOR2_X4 U2310 ( .A1(n451), .A2(n454), .ZN(n1556) );
  NAND2_X4 U2311 ( .A1(n451), .A2(n454), .ZN(n1557) );
  XOR2_X2 U2312 ( .A(n1565), .B(n1418), .Z(n2855) );
  AOI21_X4 U2313 ( .B1(n1599), .B2(n1559), .A(n1560), .ZN(n1558) );
  NOR2_X4 U2314 ( .A1(n1568), .A2(n1561), .ZN(n1559) );
  OAI21_X4 U2315 ( .B1(n1569), .B2(n1561), .A(n1564), .ZN(n1560) );
  NAND2_X4 U2318 ( .A1(n1700), .A2(n1564), .ZN(n1418) );
  NOR2_X4 U2320 ( .A1(n448), .A2(n451), .ZN(n1561) );
  NAND2_X4 U2321 ( .A1(n448), .A2(n451), .ZN(n1564) );
  XOR2_X2 U2322 ( .A(n1578), .B(n1419), .Z(n2856) );
  AOI21_X4 U2323 ( .B1(n1599), .B2(n1570), .A(n1571), .ZN(n1565) );
  NAND2_X4 U2330 ( .A1(n1586), .A2(n1574), .ZN(n1568) );
  AOI21_X4 U2331 ( .B1(n1574), .B2(n1587), .A(n1575), .ZN(n1569) );
  NOR2_X4 U2332 ( .A1(n1581), .A2(n1576), .ZN(n1574) );
  OAI21_X4 U2333 ( .B1(n1576), .B2(n1584), .A(n1577), .ZN(n1575) );
  NAND2_X4 U2334 ( .A1(n1701), .A2(n1577), .ZN(n1419) );
  NOR2_X4 U2336 ( .A1(n445), .A2(n448), .ZN(n1576) );
  NAND2_X4 U2337 ( .A1(n445), .A2(n448), .ZN(n1577) );
  XOR2_X2 U2338 ( .A(n1585), .B(n1420), .Z(n2857) );
  AOI21_X4 U2339 ( .B1(n1599), .B2(n1579), .A(n1580), .ZN(n1578) );
  NOR2_X4 U2340 ( .A1(n1588), .A2(n1581), .ZN(n1579) );
  OAI21_X4 U2341 ( .B1(n1589), .B2(n1581), .A(n1584), .ZN(n1580) );
  NAND2_X4 U2344 ( .A1(n1702), .A2(n1584), .ZN(n1420) );
  NOR2_X4 U2346 ( .A1(n442), .A2(n445), .ZN(n1581) );
  NAND2_X4 U2347 ( .A1(n442), .A2(n445), .ZN(n1584) );
  XOR2_X2 U2348 ( .A(n1594), .B(n1421), .Z(n2858) );
  AOI21_X4 U2349 ( .B1(n1599), .B2(n1586), .A(n1587), .ZN(n1585) );
  NOR2_X4 U2354 ( .A1(n1597), .A2(n1592), .ZN(n1586) );
  OAI21_X4 U2355 ( .B1(n1592), .B2(n1598), .A(n1593), .ZN(n1587) );
  NAND2_X4 U2356 ( .A1(n1703), .A2(n1593), .ZN(n1421) );
  NOR2_X4 U2358 ( .A1(n439), .A2(n442), .ZN(n1592) );
  NAND2_X4 U2359 ( .A1(n439), .A2(n442), .ZN(n1593) );
  XNOR2_X2 U2360 ( .A(n1599), .B(n1422), .ZN(n2859) );
  AOI21_X4 U2361 ( .B1(n1599), .B2(n1704), .A(n1596), .ZN(n1594) );
  NAND2_X4 U2364 ( .A1(n1704), .A2(n1598), .ZN(n1422) );
  NOR2_X4 U2366 ( .A1(n436), .A2(n439), .ZN(n1597) );
  NAND2_X4 U2367 ( .A1(n436), .A2(n439), .ZN(n1598) );
  XOR2_X2 U2368 ( .A(n1609), .B(n1423), .Z(n2860) );
  AOI21_X4 U2370 ( .B1(n1655), .B2(n1601), .A(n1602), .ZN(n1600) );
  NOR2_X4 U2371 ( .A1(n1629), .A2(n1603), .ZN(n1601) );
  OAI21_X4 U2372 ( .B1(n1630), .B2(n1603), .A(n1604), .ZN(n1602) );
  NAND2_X4 U2373 ( .A1(n1617), .A2(n1605), .ZN(n1603) );
  AOI21_X4 U2374 ( .B1(n1605), .B2(n1620), .A(n1606), .ZN(n1604) );
  NOR2_X4 U2375 ( .A1(n1612), .A2(n1607), .ZN(n1605) );
  OAI21_X4 U2376 ( .B1(n1607), .B2(n1613), .A(n1608), .ZN(n1606) );
  NAND2_X4 U2377 ( .A1(n1705), .A2(n1608), .ZN(n1423) );
  NOR2_X4 U2379 ( .A1(n433), .A2(n436), .ZN(n1607) );
  NAND2_X4 U2380 ( .A1(n433), .A2(n436), .ZN(n1608) );
  XNOR2_X2 U2381 ( .A(n1614), .B(n1424), .ZN(n2861) );
  AOI21_X4 U2382 ( .B1(n1614), .B2(n1706), .A(n1611), .ZN(n1609) );
  NAND2_X4 U2385 ( .A1(n1706), .A2(n1613), .ZN(n1424) );
  NOR2_X4 U2387 ( .A1(n430), .A2(n433), .ZN(n1612) );
  NAND2_X4 U2388 ( .A1(n430), .A2(n433), .ZN(n1613) );
  XOR2_X2 U2389 ( .A(n1623), .B(n1425), .Z(n2862) );
  OAI21_X4 U2390 ( .B1(n1654), .B2(n1615), .A(n1616), .ZN(n1614) );
  NAND2_X4 U2391 ( .A1(n1631), .A2(n1617), .ZN(n1615) );
  AOI21_X4 U2392 ( .B1(n1632), .B2(n1617), .A(n1620), .ZN(n1616) );
  NOR2_X4 U2395 ( .A1(n1626), .A2(n1621), .ZN(n1617) );
  OAI21_X4 U2396 ( .B1(n1621), .B2(n1627), .A(n1622), .ZN(n1620) );
  NAND2_X4 U2397 ( .A1(n1707), .A2(n1622), .ZN(n1425) );
  NOR2_X4 U2399 ( .A1(n427), .A2(n430), .ZN(n1621) );
  NAND2_X4 U2400 ( .A1(n427), .A2(n430), .ZN(n1622) );
  XNOR2_X2 U2401 ( .A(n1628), .B(n1426), .ZN(n2863) );
  AOI21_X4 U2402 ( .B1(n1628), .B2(n1708), .A(n1625), .ZN(n1623) );
  NAND2_X4 U2405 ( .A1(n1708), .A2(n1627), .ZN(n1426) );
  NOR2_X4 U2407 ( .A1(n424), .A2(n427), .ZN(n1626) );
  NAND2_X4 U2408 ( .A1(n424), .A2(n427), .ZN(n1627) );
  XOR2_X2 U2409 ( .A(n1639), .B(n1427), .Z(n2864) );
  OAI21_X4 U2410 ( .B1(n1654), .B2(n1629), .A(n1630), .ZN(n1628) );
  NAND2_X4 U2415 ( .A1(n1647), .A2(n1635), .ZN(n1629) );
  AOI21_X4 U2416 ( .B1(n1635), .B2(n1648), .A(n1636), .ZN(n1630) );
  NOR2_X4 U2417 ( .A1(n1642), .A2(n1637), .ZN(n1635) );
  OAI21_X4 U2418 ( .B1(n1637), .B2(n1643), .A(n1638), .ZN(n1636) );
  NAND2_X4 U2419 ( .A1(n1709), .A2(n1638), .ZN(n1427) );
  NOR2_X4 U2421 ( .A1(n421), .A2(n424), .ZN(n1637) );
  NAND2_X4 U2422 ( .A1(n421), .A2(n424), .ZN(n1638) );
  XNOR2_X2 U2423 ( .A(n1644), .B(n1428), .ZN(n2865) );
  AOI21_X4 U2424 ( .B1(n1644), .B2(n1710), .A(n1641), .ZN(n1639) );
  NAND2_X4 U2427 ( .A1(n1710), .A2(n1643), .ZN(n1428) );
  NOR2_X4 U2429 ( .A1(n418), .A2(n421), .ZN(n1642) );
  NAND2_X4 U2430 ( .A1(n418), .A2(n421), .ZN(n1643) );
  XNOR2_X2 U2431 ( .A(n1651), .B(n1429), .ZN(n2866) );
  OAI21_X4 U2432 ( .B1(n1654), .B2(n1645), .A(n1646), .ZN(n1644) );
  NOR2_X4 U2435 ( .A1(n1652), .A2(n1649), .ZN(n1647) );
  OAI21_X4 U2436 ( .B1(n1649), .B2(n1653), .A(n1650), .ZN(n1648) );
  NAND2_X4 U2437 ( .A1(n1711), .A2(n1650), .ZN(n1429) );
  NOR2_X4 U2439 ( .A1(n415), .A2(n418), .ZN(n1649) );
  NAND2_X4 U2440 ( .A1(n415), .A2(n418), .ZN(n1650) );
  XOR2_X2 U2441 ( .A(n1654), .B(n1430), .Z(n2867) );
  OAI21_X4 U2442 ( .B1(n1654), .B2(n1652), .A(n1653), .ZN(n1651) );
  NAND2_X4 U2443 ( .A1(n1712), .A2(n1653), .ZN(n1430) );
  NOR2_X4 U2445 ( .A1(n412), .A2(n415), .ZN(n1652) );
  NAND2_X4 U2446 ( .A1(n412), .A2(n415), .ZN(n1653) );
  XNOR2_X2 U2447 ( .A(n1662), .B(n1431), .ZN(n2868) );
  OAI21_X4 U2449 ( .B1(n1676), .B2(n1656), .A(n1657), .ZN(n1655) );
  NAND2_X4 U2450 ( .A1(n1666), .A2(n1658), .ZN(n1656) );
  AOI21_X4 U2451 ( .B1(n1658), .B2(n1667), .A(n1659), .ZN(n1657) );
  NOR2_X4 U2452 ( .A1(n1663), .A2(n1660), .ZN(n1658) );
  OAI21_X4 U2453 ( .B1(n1660), .B2(n1664), .A(n1661), .ZN(n1659) );
  NAND2_X4 U2454 ( .A1(n1713), .A2(n1661), .ZN(n1431) );
  NOR2_X4 U2456 ( .A1(n409), .A2(n412), .ZN(n1660) );
  NAND2_X4 U2457 ( .A1(n409), .A2(n412), .ZN(n1661) );
  XOR2_X2 U2458 ( .A(n1665), .B(n1432), .Z(n2869) );
  OAI21_X4 U2459 ( .B1(n1665), .B2(n1663), .A(n1664), .ZN(n1662) );
  NAND2_X4 U2460 ( .A1(n1714), .A2(n1664), .ZN(n1432) );
  NOR2_X4 U2462 ( .A1(n406), .A2(n409), .ZN(n1663) );
  NAND2_X4 U2463 ( .A1(n406), .A2(n409), .ZN(n1664) );
  XOR2_X2 U2464 ( .A(n1670), .B(n1433), .Z(n2870) );
  AOI21_X4 U2465 ( .B1(n1675), .B2(n1666), .A(n1667), .ZN(n1665) );
  NOR2_X4 U2466 ( .A1(n1673), .A2(n1668), .ZN(n1666) );
  OAI21_X4 U2467 ( .B1(n1668), .B2(n1674), .A(n1669), .ZN(n1667) );
  NAND2_X4 U2468 ( .A1(n1715), .A2(n1669), .ZN(n1433) );
  NOR2_X4 U2470 ( .A1(n403), .A2(n406), .ZN(n1668) );
  NAND2_X4 U2471 ( .A1(n403), .A2(n406), .ZN(n1669) );
  XNOR2_X2 U2472 ( .A(n1675), .B(n1434), .ZN(n2871) );
  AOI21_X4 U2473 ( .B1(n1675), .B2(n1716), .A(n1672), .ZN(n1670) );
  NAND2_X4 U2476 ( .A1(n1716), .A2(n1674), .ZN(n1434) );
  NOR2_X4 U2478 ( .A1(n400), .A2(n403), .ZN(n1673) );
  NAND2_X4 U2479 ( .A1(n400), .A2(n403), .ZN(n1674) );
  XNOR2_X2 U2480 ( .A(n1681), .B(n1435), .ZN(n2872) );
  AOI21_X4 U2482 ( .B1(n1677), .B2(n1685), .A(n1678), .ZN(n1676) );
  NOR2_X4 U2483 ( .A1(n1682), .A2(n1679), .ZN(n1677) );
  OAI21_X4 U2484 ( .B1(n1679), .B2(n1683), .A(n1680), .ZN(n1678) );
  NAND2_X4 U2485 ( .A1(n1717), .A2(n1680), .ZN(n1435) );
  NOR2_X4 U2487 ( .A1(n397), .A2(n400), .ZN(n1679) );
  NAND2_X4 U2488 ( .A1(n397), .A2(n400), .ZN(n1680) );
  XOR2_X2 U2489 ( .A(n1436), .B(n1684), .Z(n2873) );
  OAI21_X4 U2490 ( .B1(n1682), .B2(n1684), .A(n1683), .ZN(n1681) );
  NAND2_X4 U2491 ( .A1(n1718), .A2(n1683), .ZN(n1436) );
  NOR2_X4 U2493 ( .A1(n393), .A2(n397), .ZN(n1682) );
  NAND2_X4 U2494 ( .A1(n393), .A2(n397), .ZN(n1683) );
  NAND2_X4 U2498 ( .A1(n1719), .A2(n1684), .ZN(n2840) );
  NOR2_X4 U2500 ( .A1(n390), .A2(n393), .ZN(n1686) );
  NAND2_X4 U2501 ( .A1(n390), .A2(n393), .ZN(n1684) );
  INV_X1 U2506 ( .A(n268), .ZN(n3229) );
  INV_X1 U2507 ( .A(n265), .ZN(n3232) );
  INV_X1 U2508 ( .A(n271), .ZN(n3224) );
  XOR2_X1 U2509 ( .A(a[22]), .B(n283), .Z(n2933) );
  XNOR2_X1 U2510 ( .A(n280), .B(a[21]), .ZN(n2911) );
  XNOR2_X1 U2511 ( .A(a[21]), .B(a[22]), .ZN(n2922) );
  XOR2_X1 U2512 ( .A(a[16]), .B(n277), .Z(n2935) );
  XNOR2_X1 U2513 ( .A(a[18]), .B(a[19]), .ZN(n2923) );
  XOR2_X1 U2514 ( .A(a[1]), .B(n262), .Z(n2940) );
  XOR2_X1 U2515 ( .A(a[13]), .B(n274), .Z(n2936) );
  XNOR2_X1 U2516 ( .A(n274), .B(a[15]), .ZN(n2913) );
  XNOR2_X1 U2517 ( .A(a[15]), .B(a[16]), .ZN(n2924) );
  XNOR2_X1 U2518 ( .A(n262), .B(a[3]), .ZN(n2917) );
  INV_X1 U2519 ( .A(a[10]), .ZN(n3227) );
  XNOR2_X1 U2520 ( .A(n271), .B(a[12]), .ZN(n2914) );
  XNOR2_X1 U2521 ( .A(a[12]), .B(a[13]), .ZN(n2925) );
  XNOR2_X1 U2522 ( .A(a[3]), .B(a[4]), .ZN(n2928) );
  XNOR2_X1 U2523 ( .A(n268), .B(a[9]), .ZN(n2915) );
  XNOR2_X1 U2524 ( .A(a[9]), .B(a[10]), .ZN(n2926) );
  XOR2_X1 U2525 ( .A(a[28]), .B(n289), .Z(n2931) );
  XNOR2_X1 U2526 ( .A(n265), .B(a[6]), .ZN(n2916) );
  XNOR2_X1 U2527 ( .A(a[27]), .B(a[28]), .ZN(n2920) );
  XOR2_X1 U2528 ( .A(a[25]), .B(n286), .Z(n2932) );
  XNOR2_X1 U2529 ( .A(a[24]), .B(a[25]), .ZN(n2921) );
  INV_X1 U2530 ( .A(a[7]), .ZN(n3230) );
  XNOR2_X1 U2531 ( .A(a[6]), .B(a[7]), .ZN(n2927) );
  XNOR2_X1 U2532 ( .A(a[30]), .B(a[31]), .ZN(n2919) );
  XNOR2_X1 U2533 ( .A(a[0]), .B(a[1]), .ZN(n2929) );
  OR2_X1 U2534 ( .A1(n2929), .A2(a[0]), .ZN(n3245) );
  INV_X1 U2535 ( .A(a[0]), .ZN(n2918) );
  BUF_X1 U2536 ( .A(n336), .Z(n3126) );
  BUF_X1 U2537 ( .A(n339), .Z(n3127) );
  INV_X1 U2538 ( .A(n2917), .ZN(n3244) );
  BUF_X1 U2539 ( .A(n348), .Z(n3128) );
  BUF_X1 U2540 ( .A(n351), .Z(n3129) );
  BUF_X1 U2541 ( .A(n354), .Z(n3130) );
  XOR2_X1 U2542 ( .A(a[19]), .B(n280), .Z(n2934) );
  OR2_X1 U2543 ( .A1(n2936), .A2(n2914), .ZN(n3131) );
  INV_X1 U2544 ( .A(n3131), .ZN(n3132) );
  INV_X1 U2545 ( .A(n3131), .ZN(n3133) );
  OR2_X1 U2546 ( .A1(n2935), .A2(n2913), .ZN(n3134) );
  INV_X1 U2547 ( .A(n3134), .ZN(n3135) );
  INV_X1 U2548 ( .A(n3134), .ZN(n3136) );
  NOR2_X4 U2549 ( .A1(n2934), .A2(n2912), .ZN(n3137) );
  XNOR2_X1 U2550 ( .A(n277), .B(a[18]), .ZN(n2912) );
  NOR2_X1 U2551 ( .A1(n2934), .A2(n2912), .ZN(n303) );
  OR2_X1 U2552 ( .A1(n2933), .A2(n2911), .ZN(n3138) );
  INV_X1 U2553 ( .A(n3138), .ZN(n3139) );
  INV_X1 U2554 ( .A(n3138), .ZN(n3140) );
  OR2_X1 U2555 ( .A1(n2932), .A2(n2910), .ZN(n3141) );
  INV_X1 U2556 ( .A(n3141), .ZN(n3142) );
  INV_X1 U2557 ( .A(n3141), .ZN(n3143) );
  XNOR2_X1 U2558 ( .A(n283), .B(a[24]), .ZN(n2910) );
  OR2_X1 U2559 ( .A1(n2931), .A2(n2909), .ZN(n3144) );
  INV_X1 U2560 ( .A(n3144), .ZN(n3145) );
  INV_X1 U2561 ( .A(n3144), .ZN(n3146) );
  XNOR2_X1 U2562 ( .A(n286), .B(a[27]), .ZN(n2909) );
  OR2_X1 U2563 ( .A1(n2908), .A2(a[31]), .ZN(n3147) );
  INV_X1 U2564 ( .A(n3147), .ZN(n3148) );
  INV_X1 U2565 ( .A(n3147), .ZN(n3149) );
  XNOR2_X1 U2566 ( .A(n289), .B(a[30]), .ZN(n2908) );
  BUF_X1 U2567 ( .A(n357), .Z(n3150) );
  NAND2_X4 U2568 ( .A1(n2933), .A2(n3238), .ZN(n357) );
  AND2_X1 U2569 ( .A1(n2932), .A2(n3237), .ZN(n3151) );
  INV_X1 U2570 ( .A(n3151), .ZN(n3152) );
  INV_X4 U2571 ( .A(n3151), .ZN(n3153) );
  AND2_X1 U2572 ( .A1(n2931), .A2(n3236), .ZN(n3154) );
  INV_X1 U2573 ( .A(n3154), .ZN(n3155) );
  INV_X4 U2574 ( .A(n3154), .ZN(n3156) );
  AND2_X1 U2575 ( .A1(a[31]), .A2(n3235), .ZN(n3157) );
  INV_X1 U2576 ( .A(n3157), .ZN(n3158) );
  INV_X4 U2577 ( .A(n3157), .ZN(n3159) );
  XOR2_X1 U2578 ( .A(n719), .B(n718), .Z(n3160) );
  XOR2_X1 U2579 ( .A(n520), .B(n3160), .Z(product[62]) );
  NAND2_X1 U2580 ( .A1(n520), .A2(n719), .ZN(n3161) );
  NAND2_X1 U2581 ( .A1(n520), .A2(n718), .ZN(n3162) );
  NAND2_X1 U2582 ( .A1(n719), .A2(n718), .ZN(n3163) );
  NAND3_X1 U2583 ( .A1(n3161), .A2(n3163), .A3(n3162), .ZN(n519) );
  BUF_X1 U2584 ( .A(n536), .Z(n3164) );
  XOR2_X1 U2585 ( .A(n864), .B(n877), .Z(n3165) );
  XOR2_X1 U2586 ( .A(n539), .B(n3165), .Z(product[43]) );
  NAND2_X1 U2587 ( .A1(n539), .A2(n864), .ZN(n3166) );
  NAND2_X1 U2588 ( .A1(n539), .A2(n877), .ZN(n3167) );
  NAND2_X1 U2589 ( .A1(n864), .A2(n877), .ZN(n3168) );
  NAND3_X1 U2590 ( .A1(n3166), .A2(n3168), .A3(n3167), .ZN(n538) );
  BUF_X1 U2591 ( .A(n527), .Z(n3169) );
  BUF_X1 U2592 ( .A(n537), .Z(n3170) );
  BUF_X1 U2593 ( .A(n587), .Z(n3171) );
  BUF_X1 U2594 ( .A(n659), .Z(n3172) );
  INV_X1 U2595 ( .A(n717), .ZN(n718) );
  NAND3_X1 U2596 ( .A1(n3198), .A2(n3200), .A3(n3199), .ZN(n536) );
  AOI21_X2 U2597 ( .B1(n555), .B2(n684), .A(n552), .ZN(n550) );
  OAI21_X1 U2598 ( .B1(n660), .B2(n662), .A(n661), .ZN(n659) );
  OAI21_X2 U2599 ( .B1(n644), .B2(n646), .A(n645), .ZN(n643) );
  XNOR2_X1 U2600 ( .A(n3171), .B(n495), .ZN(product[25]) );
  XOR2_X1 U2601 ( .A(n590), .B(n496), .Z(product[24]) );
  OAI21_X2 U2602 ( .B1(n590), .B2(n588), .A(n589), .ZN(n587) );
  XNOR2_X1 U2603 ( .A(n603), .B(n499), .ZN(product[21]) );
  XNOR2_X1 U2604 ( .A(n595), .B(n497), .ZN(product[23]) );
  OAI21_X2 U2605 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  XOR2_X1 U2606 ( .A(n598), .B(n498), .Z(product[22]) );
  OAI21_X2 U2607 ( .B1(n606), .B2(n604), .A(n605), .ZN(n603) );
  BUF_X1 U2608 ( .A(n526), .Z(n3173) );
  NAND2_X1 U2609 ( .A1(n519), .A2(n3234), .ZN(n3176) );
  NAND2_X1 U2610 ( .A1(n3174), .A2(n3175), .ZN(n3177) );
  NAND2_X1 U2611 ( .A1(n3176), .A2(n3177), .ZN(product[63]) );
  INV_X1 U2612 ( .A(n519), .ZN(n3174) );
  INV_X1 U2613 ( .A(n3234), .ZN(n3175) );
  XOR2_X1 U2614 ( .A(n750), .B(n757), .Z(n3178) );
  XOR2_X1 U2615 ( .A(n528), .B(n3178), .Z(product[54]) );
  NAND2_X1 U2616 ( .A1(n528), .A2(n750), .ZN(n3179) );
  NAND2_X1 U2617 ( .A1(n528), .A2(n757), .ZN(n3180) );
  NAND2_X1 U2618 ( .A1(n750), .A2(n757), .ZN(n3181) );
  NAND3_X1 U2619 ( .A1(n3179), .A2(n3181), .A3(n3180), .ZN(n527) );
  XOR2_X1 U2620 ( .A(n851), .B(n863), .Z(n3182) );
  XOR2_X1 U2621 ( .A(n538), .B(n3182), .Z(product[44]) );
  NAND2_X1 U2622 ( .A1(n538), .A2(n851), .ZN(n3183) );
  NAND2_X1 U2623 ( .A1(n538), .A2(n863), .ZN(n3184) );
  NAND2_X1 U2624 ( .A1(n851), .A2(n863), .ZN(n3185) );
  NAND3_X1 U2625 ( .A1(n3183), .A2(n3185), .A3(n3184), .ZN(n537) );
  NAND3_X1 U2626 ( .A1(n3206), .A2(n3207), .A3(n3208), .ZN(n3186) );
  NAND3_X1 U2627 ( .A1(n3214), .A2(n3215), .A3(n3216), .ZN(n3187) );
  AOI21_X1 U2628 ( .B1(n3190), .B2(n684), .A(n552), .ZN(n3188) );
  BUF_X1 U2629 ( .A(n643), .Z(n3189) );
  BUF_X1 U2630 ( .A(n555), .Z(n3190) );
  NAND3_X1 U2631 ( .A1(n3194), .A2(n3196), .A3(n3195), .ZN(n526) );
  INV_X1 U2632 ( .A(n485), .ZN(n3234) );
  BUF_X1 U2633 ( .A(n525), .Z(n3191) );
  BUF_X1 U2634 ( .A(n535), .Z(n3192) );
  XOR2_X1 U2635 ( .A(n744), .B(n749), .Z(n3193) );
  XOR2_X1 U2636 ( .A(n3169), .B(n3193), .Z(product[55]) );
  NAND2_X1 U2637 ( .A1(n527), .A2(n744), .ZN(n3194) );
  NAND2_X1 U2638 ( .A1(n527), .A2(n749), .ZN(n3195) );
  NAND2_X1 U2639 ( .A1(n744), .A2(n749), .ZN(n3196) );
  XOR2_X1 U2640 ( .A(n837), .B(n850), .Z(n3197) );
  XOR2_X1 U2641 ( .A(n3170), .B(n3197), .Z(product[45]) );
  NAND2_X1 U2642 ( .A1(n537), .A2(n837), .ZN(n3198) );
  NAND2_X1 U2643 ( .A1(n537), .A2(n850), .ZN(n3199) );
  NAND2_X1 U2644 ( .A1(n837), .A2(n850), .ZN(n3200) );
  BUF_X1 U2645 ( .A(n3190), .Z(n3201) );
  OR2_X1 U2646 ( .A1(n2841), .A2(n342), .ZN(n3202) );
  NAND2_X1 U2647 ( .A1(n3202), .A2(n2671), .ZN(n2637) );
  BUF_X1 U2648 ( .A(n571), .Z(n3203) );
  BUF_X1 U2649 ( .A(n611), .Z(n3204) );
  NAND3_X1 U2650 ( .A1(n3206), .A2(n3207), .A3(n3208), .ZN(n525) );
  NAND3_X1 U2651 ( .A1(n3214), .A2(n3215), .A3(n3216), .ZN(n535) );
  OAI21_X1 U2652 ( .B1(n558), .B2(n556), .A(n557), .ZN(n555) );
  INV_X8 U2653 ( .A(n390), .ZN(n2841) );
  INV_X1 U2654 ( .A(n1400), .ZN(n2671) );
  OAI21_X1 U2655 ( .B1(n2839), .B2(n342), .A(n2669), .ZN(n2635) );
  AOI222_X1 U2656 ( .A1(n295), .A2(n397), .B1(n317), .B2(n393), .C1(n372), 
        .C2(n390), .ZN(n2669) );
  XOR2_X1 U2657 ( .A(n2636), .B(n268), .Z(n2022) );
  XOR2_X1 U2658 ( .A(n743), .B(n739), .Z(n3205) );
  XOR2_X1 U2659 ( .A(n3205), .B(n3173), .Z(product[56]) );
  NAND2_X2 U2660 ( .A1(n743), .A2(n739), .ZN(n3206) );
  NAND2_X1 U2661 ( .A1(n526), .A2(n743), .ZN(n3207) );
  NAND2_X1 U2662 ( .A1(n739), .A2(n526), .ZN(n3208) );
  XOR2_X1 U2663 ( .A(n738), .B(n733), .Z(n3209) );
  XOR2_X1 U2664 ( .A(n3209), .B(n3191), .Z(product[57]) );
  NAND2_X1 U2665 ( .A1(n738), .A2(n733), .ZN(n3210) );
  NAND2_X1 U2666 ( .A1(n738), .A2(n3186), .ZN(n3211) );
  NAND2_X1 U2667 ( .A1(n733), .A2(n525), .ZN(n3212) );
  NAND3_X1 U2668 ( .A1(n3210), .A2(n3211), .A3(n3212), .ZN(n524) );
  XOR2_X1 U2669 ( .A(n825), .B(n836), .Z(n3213) );
  XOR2_X1 U2670 ( .A(n3213), .B(n3164), .Z(product[46]) );
  NAND2_X2 U2671 ( .A1(n825), .A2(n836), .ZN(n3214) );
  NAND2_X1 U2672 ( .A1(n825), .A2(n536), .ZN(n3215) );
  NAND2_X1 U2673 ( .A1(n836), .A2(n536), .ZN(n3216) );
  XOR2_X1 U2674 ( .A(n814), .B(n824), .Z(n3217) );
  XOR2_X1 U2675 ( .A(n3217), .B(n3192), .Z(product[47]) );
  NAND2_X1 U2676 ( .A1(n814), .A2(n824), .ZN(n3218) );
  NAND2_X1 U2677 ( .A1(n814), .A2(n3187), .ZN(n3219) );
  NAND2_X1 U2678 ( .A1(n824), .A2(n535), .ZN(n3220) );
  NAND3_X1 U2679 ( .A1(n3218), .A2(n3219), .A3(n3220), .ZN(n534) );
  BUF_X1 U2680 ( .A(n563), .Z(n3221) );
  BUF_X1 U2681 ( .A(n579), .Z(n3222) );
  BUF_X1 U2682 ( .A(n619), .Z(n3223) );
  OAI21_X1 U2683 ( .B1(n2840), .B2(n342), .A(n2670), .ZN(n2636) );
  AOI22_X1 U2684 ( .A1(n295), .A2(n393), .B1(n317), .B2(n390), .ZN(n2670) );
  XNOR2_X1 U2685 ( .A(n2569), .B(n3224), .ZN(n1988) );
  INV_X2 U2686 ( .A(n291), .ZN(n3225) );
  INV_X8 U2687 ( .A(n3225), .ZN(n3226) );
  NOR2_X1 U2688 ( .A1(n2940), .A2(n2918), .ZN(n291) );
  NAND2_X4 U2689 ( .A1(n2934), .A2(n3239), .ZN(n354) );
  INV_X8 U2690 ( .A(n3248), .ZN(n319) );
  NOR2_X1 U2691 ( .A1(n1339), .A2(n1344), .ZN(n641) );
  NAND2_X2 U2692 ( .A1(n1339), .A2(n1344), .ZN(n642) );
  OAI21_X1 U2693 ( .B1(n2841), .B2(n345), .A(n2603), .ZN(n2569) );
  XNOR2_X2 U2694 ( .A(n3227), .B(n271), .ZN(n2937) );
  OR2_X4 U2695 ( .A1(n2939), .A2(n2917), .ZN(n3228) );
  INV_X32 U2696 ( .A(n3228), .ZN(n293) );
  XNOR2_X1 U2697 ( .A(n2637), .B(n3229), .ZN(n2023) );
  NOR2_X2 U2698 ( .A1(n1373), .A2(n2090), .ZN(n673) );
  NAND2_X2 U2699 ( .A1(n1373), .A2(n2090), .ZN(n674) );
  XNOR2_X2 U2700 ( .A(n3230), .B(n268), .ZN(n2938) );
  NOR2_X1 U2701 ( .A1(n1351), .A2(n1356), .ZN(n649) );
  NAND2_X2 U2702 ( .A1(n1351), .A2(n1356), .ZN(n650) );
  INV_X8 U2703 ( .A(n3246), .ZN(n315) );
  OR2_X4 U2704 ( .A1(n2937), .A2(n2915), .ZN(n3231) );
  INV_X32 U2705 ( .A(n3231), .ZN(n297) );
  INV_X8 U2706 ( .A(n3247), .ZN(n317) );
  XNOR2_X2 U2707 ( .A(n2705), .B(n3232), .ZN(n2058) );
  NAND2_X4 U2708 ( .A1(n2935), .A2(n3240), .ZN(n351) );
  XNOR2_X1 U2709 ( .A(n513), .B(n3172), .ZN(product[7]) );
  XNOR2_X1 U2710 ( .A(n651), .B(n511), .ZN(product[9]) );
  OR2_X4 U2711 ( .A1(n2938), .A2(n2916), .ZN(n3233) );
  INV_X32 U2712 ( .A(n3233), .ZN(n295) );
  XNOR2_X1 U2713 ( .A(n3221), .B(n489), .ZN(product[31]) );
  XNOR2_X1 U2714 ( .A(n3189), .B(n509), .ZN(product[11]) );
  NAND2_X4 U2715 ( .A1(n2936), .A2(n3241), .ZN(n348) );
  AOI21_X4 U2716 ( .B1(n571), .B2(n688), .A(n568), .ZN(n566) );
  XOR2_X1 U2717 ( .A(n566), .B(n490), .Z(product[30]) );
  OAI21_X2 U2718 ( .B1(n566), .B2(n564), .A(n565), .ZN(n563) );
  XOR2_X1 U2719 ( .A(n3188), .B(n486), .Z(product[34]) );
  OAI21_X1 U2720 ( .B1(n550), .B2(n548), .A(n549), .ZN(n547) );
  XOR2_X1 U2721 ( .A(n2501), .B(n274), .Z(n1953) );
  NAND2_X4 U2722 ( .A1(n2940), .A2(a[0]), .ZN(n336) );
  NAND2_X4 U2723 ( .A1(n2937), .A2(n3242), .ZN(n345) );
  XNOR2_X1 U2724 ( .A(n3203), .B(n491), .ZN(product[29]) );
  XNOR2_X1 U2725 ( .A(n3222), .B(n493), .ZN(product[27]) );
  XNOR2_X1 U2726 ( .A(n3223), .B(n503), .ZN(product[17]) );
  XNOR2_X1 U2727 ( .A(n3201), .B(n487), .ZN(product[33]) );
  XNOR2_X1 U2728 ( .A(n3204), .B(n501), .ZN(product[19]) );
  XOR2_X1 U2729 ( .A(n510), .B(n646), .Z(product[10]) );
  NAND2_X4 U2730 ( .A1(n2938), .A2(n3243), .ZN(n342) );
  NAND2_X4 U2731 ( .A1(n2939), .A2(n3244), .ZN(n339) );
  OAI21_X2 U2732 ( .B1(n654), .B2(n652), .A(n653), .ZN(n651) );
  OAI21_X2 U2733 ( .B1(n614), .B2(n612), .A(n613), .ZN(n611) );
  OAI21_X2 U2734 ( .B1(n582), .B2(n580), .A(n581), .ZN(n579) );
  OAI21_X2 U2735 ( .B1(n574), .B2(n572), .A(n573), .ZN(n571) );
  OAI21_X2 U2736 ( .B1(n622), .B2(n620), .A(n621), .ZN(n619) );
  INV_X2 U2737 ( .A(n518), .ZN(product[0]) );
  INV_X2 U2738 ( .A(n941), .ZN(n959) );
  INV_X2 U2739 ( .A(n907), .ZN(n908) );
  INV_X2 U2740 ( .A(n891), .ZN(n892) );
  INV_X2 U2741 ( .A(n848), .ZN(n862) );
  INV_X2 U2742 ( .A(n811), .ZN(n823) );
  INV_X2 U2743 ( .A(n780), .ZN(n790) );
  INV_X2 U2744 ( .A(n755), .ZN(n763) );
  INV_X2 U2745 ( .A(n736), .ZN(n742) );
  INV_X2 U2746 ( .A(n723), .ZN(n727) );
  INV_X2 U2747 ( .A(n1720), .ZN(n716) );
  INV_X2 U2748 ( .A(n681), .ZN(n715) );
  INV_X2 U2749 ( .A(n668), .ZN(n713) );
  INV_X2 U2750 ( .A(n660), .ZN(n711) );
  INV_X2 U2751 ( .A(n652), .ZN(n709) );
  INV_X2 U2752 ( .A(n644), .ZN(n707) );
  INV_X2 U2753 ( .A(n636), .ZN(n705) );
  INV_X2 U2754 ( .A(n628), .ZN(n703) );
  INV_X2 U2755 ( .A(n620), .ZN(n701) );
  INV_X2 U2756 ( .A(n612), .ZN(n699) );
  INV_X2 U2757 ( .A(n604), .ZN(n697) );
  INV_X2 U2758 ( .A(n596), .ZN(n695) );
  INV_X2 U2759 ( .A(n588), .ZN(n693) );
  INV_X2 U2760 ( .A(n580), .ZN(n691) );
  INV_X2 U2761 ( .A(n572), .ZN(n689) );
  INV_X2 U2762 ( .A(n564), .ZN(n687) );
  INV_X2 U2763 ( .A(n556), .ZN(n685) );
  INV_X2 U2764 ( .A(n548), .ZN(n683) );
  INV_X2 U2765 ( .A(n682), .ZN(n680) );
  INV_X2 U2766 ( .A(n678), .ZN(n679) );
  INV_X2 U2767 ( .A(n2091), .ZN(n676) );
  INV_X2 U2768 ( .A(n674), .ZN(n672) );
  INV_X2 U2769 ( .A(n673), .ZN(n714) );
  INV_X2 U2770 ( .A(n666), .ZN(n664) );
  INV_X2 U2771 ( .A(n665), .ZN(n712) );
  INV_X2 U2772 ( .A(n658), .ZN(n656) );
  INV_X2 U2773 ( .A(n657), .ZN(n710) );
  INV_X2 U2774 ( .A(n650), .ZN(n648) );
  INV_X2 U2775 ( .A(n649), .ZN(n708) );
  INV_X2 U2776 ( .A(n642), .ZN(n640) );
  INV_X2 U2777 ( .A(n641), .ZN(n706) );
  INV_X2 U2778 ( .A(n634), .ZN(n632) );
  INV_X2 U2779 ( .A(n633), .ZN(n704) );
  INV_X2 U2780 ( .A(n626), .ZN(n624) );
  INV_X2 U2781 ( .A(n625), .ZN(n702) );
  INV_X2 U2782 ( .A(n618), .ZN(n616) );
  INV_X2 U2783 ( .A(n617), .ZN(n700) );
  INV_X2 U2784 ( .A(n610), .ZN(n608) );
  INV_X2 U2785 ( .A(n609), .ZN(n698) );
  INV_X2 U2786 ( .A(n602), .ZN(n600) );
  INV_X2 U2787 ( .A(n601), .ZN(n696) );
  INV_X2 U2788 ( .A(n594), .ZN(n592) );
  INV_X2 U2789 ( .A(n593), .ZN(n694) );
  INV_X2 U2790 ( .A(n586), .ZN(n584) );
  INV_X2 U2791 ( .A(n585), .ZN(n692) );
  INV_X2 U2792 ( .A(n578), .ZN(n576) );
  INV_X2 U2793 ( .A(n577), .ZN(n690) );
  INV_X2 U2794 ( .A(n570), .ZN(n568) );
  INV_X2 U2795 ( .A(n569), .ZN(n688) );
  INV_X2 U2796 ( .A(n562), .ZN(n560) );
  INV_X2 U2797 ( .A(n561), .ZN(n686) );
  INV_X2 U2798 ( .A(n554), .ZN(n552) );
  INV_X2 U2799 ( .A(n553), .ZN(n684) );
  INV_X2 U2800 ( .A(n2873), .ZN(n2839) );
  INV_X2 U2801 ( .A(n2872), .ZN(n2838) );
  INV_X2 U2802 ( .A(n2871), .ZN(n2837) );
  INV_X2 U2803 ( .A(n2870), .ZN(n2836) );
  INV_X2 U2804 ( .A(n2869), .ZN(n2835) );
  INV_X2 U2805 ( .A(n2868), .ZN(n2834) );
  INV_X2 U2806 ( .A(n2867), .ZN(n2833) );
  INV_X2 U2807 ( .A(n2866), .ZN(n2832) );
  INV_X2 U2808 ( .A(n2865), .ZN(n2831) );
  INV_X2 U2809 ( .A(n2864), .ZN(n2830) );
  INV_X2 U2810 ( .A(n2863), .ZN(n2829) );
  INV_X2 U2811 ( .A(n2862), .ZN(n2828) );
  INV_X2 U2812 ( .A(n2861), .ZN(n2827) );
  INV_X2 U2813 ( .A(n2860), .ZN(n2826) );
  INV_X2 U2814 ( .A(n2859), .ZN(n2825) );
  INV_X2 U2815 ( .A(n2858), .ZN(n2824) );
  INV_X2 U2816 ( .A(n2857), .ZN(n2823) );
  INV_X2 U2817 ( .A(n2856), .ZN(n2822) );
  INV_X2 U2818 ( .A(n2855), .ZN(n2821) );
  INV_X2 U2819 ( .A(n2854), .ZN(n2820) );
  INV_X2 U2820 ( .A(n2853), .ZN(n2819) );
  INV_X2 U2821 ( .A(n2852), .ZN(n2818) );
  INV_X2 U2822 ( .A(n2851), .ZN(n2817) );
  INV_X2 U2823 ( .A(n2850), .ZN(n2816) );
  INV_X2 U2824 ( .A(n2849), .ZN(n2815) );
  INV_X2 U2825 ( .A(n2848), .ZN(n2814) );
  INV_X2 U2826 ( .A(n2847), .ZN(n2813) );
  INV_X2 U2827 ( .A(n2846), .ZN(n2812) );
  INV_X2 U2828 ( .A(n2845), .ZN(n2811) );
  INV_X2 U2829 ( .A(n2844), .ZN(n2810) );
  INV_X2 U2830 ( .A(n2843), .ZN(n2809) );
  INV_X2 U2831 ( .A(n1406), .ZN(n2807) );
  AOI22_X2 U2832 ( .A1(n3226), .A2(n393), .B1(n313), .B2(n390), .ZN(n2806) );
  INV_X2 U2833 ( .A(n3245), .ZN(n313) );
  INV_X2 U2834 ( .A(n1403), .ZN(n2739) );
  AOI22_X2 U2835 ( .A1(n293), .A2(n393), .B1(n315), .B2(n390), .ZN(n2738) );
  OR2_X2 U2836 ( .A1(n2928), .A2(n3244), .ZN(n3246) );
  OR2_X2 U2837 ( .A1(n2927), .A2(n3243), .ZN(n3247) );
  INV_X2 U2838 ( .A(n2916), .ZN(n3243) );
  INV_X2 U2839 ( .A(n1397), .ZN(n2603) );
  AOI22_X2 U2840 ( .A1(n297), .A2(n393), .B1(n319), .B2(n390), .ZN(n2602) );
  OR2_X2 U2841 ( .A1(n2926), .A2(n3242), .ZN(n3248) );
  INV_X2 U2842 ( .A(n2915), .ZN(n3242) );
  INV_X2 U2843 ( .A(n1394), .ZN(n2535) );
  AOI22_X2 U2844 ( .A1(n3133), .A2(n393), .B1(n321), .B2(n390), .ZN(n2534) );
  INV_X2 U2845 ( .A(n3249), .ZN(n321) );
  OR2_X2 U2846 ( .A1(n2925), .A2(n3241), .ZN(n3249) );
  INV_X2 U2847 ( .A(n2914), .ZN(n3241) );
  INV_X2 U2848 ( .A(n1391), .ZN(n2467) );
  AOI22_X2 U2849 ( .A1(n3136), .A2(n393), .B1(n323), .B2(n390), .ZN(n2466) );
  INV_X2 U2850 ( .A(n3250), .ZN(n323) );
  OR2_X2 U2851 ( .A1(n2924), .A2(n3240), .ZN(n3250) );
  INV_X2 U2852 ( .A(n2913), .ZN(n3240) );
  INV_X2 U2853 ( .A(n1388), .ZN(n2399) );
  AOI22_X2 U2854 ( .A1(n303), .A2(n393), .B1(n325), .B2(n390), .ZN(n2398) );
  INV_X2 U2855 ( .A(n3251), .ZN(n325) );
  OR2_X2 U2856 ( .A1(n2923), .A2(n3239), .ZN(n3251) );
  INV_X2 U2857 ( .A(n2912), .ZN(n3239) );
  INV_X2 U2858 ( .A(n1385), .ZN(n2331) );
  AOI22_X2 U2859 ( .A1(n3140), .A2(n393), .B1(n327), .B2(n390), .ZN(n2330) );
  INV_X2 U2860 ( .A(n3252), .ZN(n327) );
  OR2_X2 U2861 ( .A1(n2922), .A2(n3238), .ZN(n3252) );
  INV_X2 U2862 ( .A(n2911), .ZN(n3238) );
  INV_X2 U2863 ( .A(n1382), .ZN(n2263) );
  AOI22_X2 U2864 ( .A1(n3143), .A2(n393), .B1(n329), .B2(n390), .ZN(n2262) );
  INV_X2 U2865 ( .A(n3253), .ZN(n329) );
  OR2_X2 U2866 ( .A1(n2921), .A2(n3237), .ZN(n3253) );
  INV_X2 U2867 ( .A(n2910), .ZN(n3237) );
  INV_X2 U2868 ( .A(n1379), .ZN(n2195) );
  AOI22_X2 U2869 ( .A1(n3146), .A2(n393), .B1(n331), .B2(n390), .ZN(n2194) );
  INV_X2 U2870 ( .A(n3254), .ZN(n331) );
  OR2_X2 U2871 ( .A1(n2920), .A2(n3236), .ZN(n3254) );
  INV_X2 U2872 ( .A(n2909), .ZN(n3236) );
  INV_X2 U2873 ( .A(n1376), .ZN(n2127) );
  AOI22_X2 U2874 ( .A1(n3148), .A2(n393), .B1(n333), .B2(n390), .ZN(n2126) );
  INV_X2 U2875 ( .A(n3255), .ZN(n333) );
  OR2_X2 U2876 ( .A1(n2919), .A2(n3235), .ZN(n3255) );
  INV_X2 U2877 ( .A(n2908), .ZN(n3235) );
  INV_X2 U2878 ( .A(n262), .ZN(n2059) );
  INV_X2 U2879 ( .A(n274), .ZN(n1919) );
  INV_X2 U2880 ( .A(n277), .ZN(n1884) );
  INV_X2 U2881 ( .A(n280), .ZN(n1849) );
  INV_X2 U2882 ( .A(n283), .ZN(n1814) );
  INV_X2 U2883 ( .A(n286), .ZN(n1779) );
  INV_X2 U2884 ( .A(n289), .ZN(n1745) );
  INV_X2 U2885 ( .A(n1686), .ZN(n1719) );
  INV_X2 U2886 ( .A(n1682), .ZN(n1718) );
  INV_X2 U2887 ( .A(n1679), .ZN(n1717) );
  INV_X2 U2888 ( .A(n1668), .ZN(n1715) );
  INV_X2 U2889 ( .A(n1663), .ZN(n1714) );
  INV_X2 U2890 ( .A(n1660), .ZN(n1713) );
  INV_X2 U2891 ( .A(n1652), .ZN(n1712) );
  INV_X2 U2892 ( .A(n1649), .ZN(n1711) );
  INV_X2 U2893 ( .A(n1637), .ZN(n1709) );
  INV_X2 U2894 ( .A(n1621), .ZN(n1707) );
  INV_X2 U2895 ( .A(n1607), .ZN(n1705) );
  INV_X2 U2896 ( .A(n1592), .ZN(n1703) );
  INV_X2 U2897 ( .A(n1581), .ZN(n1702) );
  INV_X2 U2898 ( .A(n1576), .ZN(n1701) );
  INV_X2 U2899 ( .A(n1561), .ZN(n1700) );
  INV_X2 U2900 ( .A(n1556), .ZN(n1699) );
  INV_X2 U2901 ( .A(n1543), .ZN(n1698) );
  INV_X2 U2902 ( .A(n1538), .ZN(n1697) );
  INV_X2 U2903 ( .A(n1523), .ZN(n1696) );
  INV_X2 U2904 ( .A(n1518), .ZN(n1695) );
  INV_X2 U2905 ( .A(n1496), .ZN(n1693) );
  INV_X2 U2906 ( .A(n1474), .ZN(n1691) );
  INV_X2 U2907 ( .A(n1459), .ZN(n1690) );
  INV_X2 U2908 ( .A(n1450), .ZN(n1689) );
  INV_X2 U2909 ( .A(n1684), .ZN(n1685) );
  INV_X2 U2910 ( .A(n1676), .ZN(n1675) );
  INV_X2 U2911 ( .A(n1674), .ZN(n1672) );
  INV_X2 U2912 ( .A(n1673), .ZN(n1716) );
  INV_X2 U2913 ( .A(n1655), .ZN(n1654) );
  INV_X2 U2914 ( .A(n1648), .ZN(n1646) );
  INV_X2 U2915 ( .A(n1647), .ZN(n1645) );
  INV_X2 U2916 ( .A(n1643), .ZN(n1641) );
  INV_X2 U2917 ( .A(n1642), .ZN(n1710) );
  INV_X2 U2918 ( .A(n1630), .ZN(n1632) );
  INV_X2 U2919 ( .A(n1629), .ZN(n1631) );
  INV_X2 U2920 ( .A(n1627), .ZN(n1625) );
  INV_X2 U2921 ( .A(n1626), .ZN(n1708) );
  INV_X2 U2922 ( .A(n1613), .ZN(n1611) );
  INV_X2 U2923 ( .A(n1612), .ZN(n1706) );
  INV_X2 U2924 ( .A(n1600), .ZN(n1599) );
  INV_X2 U2925 ( .A(n1598), .ZN(n1596) );
  INV_X2 U2926 ( .A(n1597), .ZN(n1704) );
  INV_X2 U2927 ( .A(n1587), .ZN(n1589) );
  INV_X2 U2928 ( .A(n1586), .ZN(n1588) );
  INV_X2 U2929 ( .A(n1569), .ZN(n1571) );
  INV_X2 U2930 ( .A(n1568), .ZN(n1570) );
  INV_X2 U2931 ( .A(n1551), .ZN(n1549) );
  INV_X2 U2932 ( .A(n1550), .ZN(n1548) );
  INV_X2 U2933 ( .A(n1529), .ZN(n1531) );
  INV_X2 U2934 ( .A(n1528), .ZN(n1530) );
  INV_X2 U2935 ( .A(n1513), .ZN(n1511) );
  INV_X2 U2936 ( .A(n1512), .ZN(n1510) );
  INV_X2 U2937 ( .A(n1506), .ZN(n1504) );
  INV_X2 U2938 ( .A(n1505), .ZN(n1694) );
  INV_X2 U2939 ( .A(n1489), .ZN(n1491) );
  INV_X2 U2940 ( .A(n1488), .ZN(n1490) );
  INV_X2 U2941 ( .A(n1484), .ZN(n1482) );
  INV_X2 U2942 ( .A(n1483), .ZN(n1692) );
  INV_X2 U2943 ( .A(n1469), .ZN(n1471) );
  INV_X2 U2944 ( .A(n1468), .ZN(n1470) );
  INV_X2 U2945 ( .A(n484), .ZN(n1440) );
endmodule


module mul32_1_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n262, n265, n268, n271, n274, n277, n280, n283, n286, n289, n293,
         n295, n297, n313, n315, n317, n319, n321, n323, n325, n327, n329,
         n331, n333, n336, n339, n342, n345, n348, n351, n354, n357, n368,
         n370, n372, n374, n376, n378, n380, n382, n384, n386, n388, n390,
         n393, n397, n400, n403, n406, n409, n412, n415, n418, n421, n424,
         n427, n430, n433, n436, n439, n442, n445, n448, n451, n454, n457,
         n460, n463, n466, n469, n472, n475, n478, n481, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n552, n553,
         n554, n555, n556, n557, n558, n560, n561, n562, n563, n564, n565,
         n566, n568, n569, n570, n571, n572, n573, n574, n576, n577, n578,
         n579, n580, n581, n582, n584, n585, n586, n587, n588, n589, n590,
         n592, n593, n594, n595, n596, n597, n598, n600, n601, n602, n603,
         n604, n605, n606, n608, n609, n610, n611, n612, n613, n614, n616,
         n617, n618, n619, n620, n621, n622, n624, n625, n626, n627, n628,
         n629, n630, n632, n633, n634, n635, n636, n637, n638, n640, n641,
         n642, n643, n644, n645, n646, n648, n649, n650, n651, n652, n653,
         n654, n656, n657, n658, n659, n660, n661, n662, n664, n665, n666,
         n667, n668, n669, n670, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1376, n1377, n1379, n1380, n1382, n1383, n1385, n1386, n1388, n1389,
         n1391, n1392, n1394, n1395, n1397, n1398, n1400, n1401, n1403, n1404,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1518, n1519, n1520,
         n1521, n1522, n1523, n1526, n1527, n1528, n1529, n1530, n1531, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1564, n1565, n1568, n1569, n1570, n1571, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1584, n1585, n1586,
         n1587, n1588, n1589, n1592, n1593, n1594, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1620, n1621, n1622,
         n1623, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1635,
         n1636, n1637, n1638, n1639, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240;
  assign n262 = a[2];
  assign n265 = a[5];
  assign n268 = a[8];
  assign n271 = a[11];
  assign n274 = a[14];
  assign n277 = a[17];
  assign n280 = a[20];
  assign n283 = a[23];
  assign n286 = a[26];
  assign n289 = a[29];
  assign n390 = b[0];
  assign n393 = b[1];
  assign n397 = b[2];
  assign n400 = b[3];
  assign n403 = b[4];
  assign n406 = b[5];
  assign n409 = b[6];
  assign n412 = b[7];
  assign n415 = b[8];
  assign n418 = b[9];
  assign n421 = b[10];
  assign n424 = b[11];
  assign n427 = b[12];
  assign n430 = b[13];
  assign n433 = b[14];
  assign n436 = b[15];
  assign n439 = b[16];
  assign n442 = b[17];
  assign n445 = b[18];
  assign n448 = b[19];
  assign n451 = b[20];
  assign n454 = b[21];
  assign n457 = b[22];
  assign n460 = b[23];
  assign n463 = b[24];
  assign n466 = b[25];
  assign n469 = b[26];
  assign n472 = b[27];
  assign n475 = b[28];
  assign n478 = b[29];
  assign n481 = b[30];
  assign n484 = b[31];

  XOR2_X2 U304 ( .A(n717), .B(n716), .Z(n485) );
  FA_X1 U309 ( .A(n729), .B(n732), .CI(n524), .CO(n523), .S(product[58]) );
  FA_X1 U312 ( .A(n738), .B(n733), .CI(n525), .CO(n524), .S(product[57]) );
  FA_X1 U313 ( .A(n743), .B(n739), .CI(n526), .CO(n525), .S(product[56]) );
  FA_X1 U314 ( .A(n744), .B(n749), .CI(n527), .CO(n526), .S(product[55]) );
  FA_X1 U315 ( .A(n750), .B(n757), .CI(n528), .CO(n527), .S(product[54]) );
  FA_X1 U316 ( .A(n758), .B(n764), .CI(n529), .CO(n528), .S(product[53]) );
  FA_X1 U319 ( .A(n783), .B(n791), .CI(n532), .CO(n531), .S(product[50]) );
  FA_X1 U320 ( .A(n792), .B(n801), .CI(n533), .CO(n532), .S(product[49]) );
  FA_X1 U321 ( .A(n802), .B(n813), .CI(n534), .CO(n533), .S(product[48]) );
  FA_X1 U322 ( .A(n814), .B(n824), .CI(n535), .CO(n534), .S(product[47]) );
  FA_X1 U323 ( .A(n825), .B(n836), .CI(n536), .CO(n535), .S(product[46]) );
  FA_X1 U324 ( .A(n837), .B(n850), .CI(n537), .CO(n536), .S(product[45]) );
  FA_X1 U325 ( .A(n851), .B(n863), .CI(n538), .CO(n537), .S(product[44]) );
  FA_X1 U326 ( .A(n864), .B(n877), .CI(n539), .CO(n538), .S(product[43]) );
  FA_X1 U327 ( .A(n878), .B(n893), .CI(n540), .CO(n539), .S(product[42]) );
  FA_X1 U328 ( .A(n894), .B(n909), .CI(n541), .CO(n540), .S(product[41]) );
  FA_X1 U329 ( .A(n910), .B(n925), .CI(n542), .CO(n541), .S(product[40]) );
  FA_X1 U330 ( .A(n926), .B(n943), .CI(n543), .CO(n542), .S(product[39]) );
  NAND2_X4 U337 ( .A1(n683), .A2(n549), .ZN(n486) );
  NOR2_X4 U339 ( .A1(n1015), .A2(n1032), .ZN(n548) );
  NAND2_X4 U340 ( .A1(n1015), .A2(n1032), .ZN(n549) );
  NAND2_X4 U345 ( .A1(n684), .A2(n554), .ZN(n487) );
  NOR2_X4 U347 ( .A1(n1033), .A2(n1050), .ZN(n553) );
  NAND2_X4 U348 ( .A1(n1033), .A2(n1050), .ZN(n554) );
  NAND2_X4 U351 ( .A1(n685), .A2(n557), .ZN(n488) );
  NOR2_X4 U353 ( .A1(n1051), .A2(n1068), .ZN(n556) );
  NAND2_X4 U354 ( .A1(n1051), .A2(n1068), .ZN(n557) );
  NAND2_X4 U359 ( .A1(n686), .A2(n562), .ZN(n489) );
  NOR2_X4 U361 ( .A1(n1069), .A2(n1086), .ZN(n561) );
  NAND2_X4 U362 ( .A1(n1069), .A2(n1086), .ZN(n562) );
  NAND2_X4 U365 ( .A1(n687), .A2(n565), .ZN(n490) );
  NOR2_X4 U367 ( .A1(n1087), .A2(n1104), .ZN(n564) );
  NAND2_X4 U368 ( .A1(n1087), .A2(n1104), .ZN(n565) );
  NAND2_X4 U373 ( .A1(n688), .A2(n570), .ZN(n491) );
  NOR2_X4 U375 ( .A1(n1105), .A2(n1122), .ZN(n569) );
  NAND2_X4 U376 ( .A1(n1105), .A2(n1122), .ZN(n570) );
  NAND2_X4 U379 ( .A1(n689), .A2(n573), .ZN(n492) );
  NOR2_X4 U381 ( .A1(n1123), .A2(n1140), .ZN(n572) );
  NAND2_X4 U382 ( .A1(n1123), .A2(n1140), .ZN(n573) );
  NAND2_X4 U387 ( .A1(n690), .A2(n578), .ZN(n493) );
  NOR2_X4 U389 ( .A1(n1141), .A2(n1158), .ZN(n577) );
  NAND2_X4 U390 ( .A1(n1141), .A2(n1158), .ZN(n578) );
  NAND2_X4 U393 ( .A1(n691), .A2(n581), .ZN(n494) );
  NOR2_X4 U395 ( .A1(n1159), .A2(n1174), .ZN(n580) );
  NAND2_X4 U396 ( .A1(n1159), .A2(n1174), .ZN(n581) );
  NAND2_X4 U401 ( .A1(n692), .A2(n586), .ZN(n495) );
  NOR2_X4 U403 ( .A1(n1175), .A2(n1190), .ZN(n585) );
  NAND2_X4 U404 ( .A1(n1175), .A2(n1190), .ZN(n586) );
  XOR2_X2 U405 ( .A(n590), .B(n496), .Z(product[24]) );
  NAND2_X4 U407 ( .A1(n693), .A2(n589), .ZN(n496) );
  NOR2_X4 U409 ( .A1(n1191), .A2(n1206), .ZN(n588) );
  NAND2_X4 U412 ( .A1(n1191), .A2(n1206), .ZN(n589) );
  AOI21_X4 U414 ( .B1(n595), .B2(n694), .A(n592), .ZN(n590) );
  NAND2_X4 U417 ( .A1(n694), .A2(n594), .ZN(n497) );
  NOR2_X4 U419 ( .A1(n1207), .A2(n1220), .ZN(n593) );
  NAND2_X4 U420 ( .A1(n1207), .A2(n1220), .ZN(n594) );
  NAND2_X4 U423 ( .A1(n695), .A2(n597), .ZN(n498) );
  NOR2_X4 U425 ( .A1(n1221), .A2(n1234), .ZN(n596) );
  NAND2_X4 U426 ( .A1(n1221), .A2(n1234), .ZN(n597) );
  NAND2_X4 U431 ( .A1(n696), .A2(n602), .ZN(n499) );
  NOR2_X4 U433 ( .A1(n1235), .A2(n1248), .ZN(n601) );
  NAND2_X4 U434 ( .A1(n1235), .A2(n1248), .ZN(n602) );
  XOR2_X2 U435 ( .A(n606), .B(n500), .Z(product[20]) );
  NAND2_X4 U437 ( .A1(n697), .A2(n605), .ZN(n500) );
  NOR2_X4 U439 ( .A1(n1249), .A2(n1260), .ZN(n604) );
  NAND2_X4 U440 ( .A1(n1249), .A2(n1260), .ZN(n605) );
  AOI21_X4 U442 ( .B1(n611), .B2(n698), .A(n608), .ZN(n606) );
  NAND2_X4 U445 ( .A1(n698), .A2(n610), .ZN(n501) );
  NOR2_X4 U447 ( .A1(n1261), .A2(n1272), .ZN(n609) );
  NAND2_X4 U448 ( .A1(n1261), .A2(n1272), .ZN(n610) );
  NAND2_X4 U451 ( .A1(n699), .A2(n613), .ZN(n502) );
  NOR2_X4 U453 ( .A1(n1273), .A2(n1284), .ZN(n612) );
  NAND2_X4 U454 ( .A1(n1273), .A2(n1284), .ZN(n613) );
  AOI21_X4 U456 ( .B1(n619), .B2(n700), .A(n616), .ZN(n614) );
  NAND2_X4 U459 ( .A1(n700), .A2(n618), .ZN(n503) );
  NOR2_X4 U461 ( .A1(n1285), .A2(n1294), .ZN(n617) );
  NAND2_X4 U462 ( .A1(n1285), .A2(n1294), .ZN(n618) );
  NAND2_X4 U465 ( .A1(n701), .A2(n621), .ZN(n504) );
  NOR2_X4 U467 ( .A1(n1295), .A2(n1304), .ZN(n620) );
  NAND2_X4 U468 ( .A1(n1295), .A2(n1304), .ZN(n621) );
  NAND2_X4 U473 ( .A1(n702), .A2(n626), .ZN(n505) );
  NOR2_X4 U475 ( .A1(n1305), .A2(n1314), .ZN(n625) );
  NAND2_X4 U476 ( .A1(n1305), .A2(n1314), .ZN(n626) );
  NAND2_X4 U479 ( .A1(n703), .A2(n629), .ZN(n506) );
  NOR2_X4 U481 ( .A1(n1315), .A2(n1322), .ZN(n628) );
  NAND2_X4 U482 ( .A1(n1315), .A2(n1322), .ZN(n629) );
  NAND2_X4 U487 ( .A1(n704), .A2(n634), .ZN(n507) );
  NOR2_X4 U489 ( .A1(n1323), .A2(n1330), .ZN(n633) );
  NAND2_X4 U490 ( .A1(n1323), .A2(n1330), .ZN(n634) );
  NAND2_X4 U493 ( .A1(n705), .A2(n637), .ZN(n508) );
  NOR2_X4 U495 ( .A1(n1331), .A2(n1338), .ZN(n636) );
  NAND2_X4 U496 ( .A1(n1331), .A2(n1338), .ZN(n637) );
  NAND2_X4 U501 ( .A1(n706), .A2(n642), .ZN(n509) );
  NAND2_X4 U504 ( .A1(n1339), .A2(n1344), .ZN(n642) );
  NAND2_X4 U507 ( .A1(n707), .A2(n645), .ZN(n510) );
  NOR2_X4 U509 ( .A1(n1345), .A2(n1350), .ZN(n644) );
  NAND2_X4 U510 ( .A1(n1345), .A2(n1350), .ZN(n645) );
  NAND2_X4 U515 ( .A1(n708), .A2(n650), .ZN(n511) );
  XOR2_X2 U519 ( .A(n654), .B(n512), .Z(product[8]) );
  NAND2_X4 U521 ( .A1(n709), .A2(n653), .ZN(n512) );
  NOR2_X4 U523 ( .A1(n1357), .A2(n1360), .ZN(n652) );
  NAND2_X4 U524 ( .A1(n1357), .A2(n1360), .ZN(n653) );
  AOI21_X4 U526 ( .B1(n659), .B2(n710), .A(n656), .ZN(n654) );
  NAND2_X4 U529 ( .A1(n710), .A2(n658), .ZN(n513) );
  NOR2_X4 U531 ( .A1(n1361), .A2(n1364), .ZN(n657) );
  NAND2_X4 U532 ( .A1(n1361), .A2(n1364), .ZN(n658) );
  XOR2_X2 U533 ( .A(n514), .B(n662), .Z(product[6]) );
  NAND2_X4 U535 ( .A1(n711), .A2(n661), .ZN(n514) );
  NAND2_X4 U538 ( .A1(n1365), .A2(n2087), .ZN(n661) );
  XNOR2_X2 U539 ( .A(n515), .B(n667), .ZN(product[5]) );
  AOI21_X4 U540 ( .B1(n712), .B2(n667), .A(n664), .ZN(n662) );
  NAND2_X4 U543 ( .A1(n712), .A2(n666), .ZN(n515) );
  NOR2_X4 U545 ( .A1(n2088), .A2(n1369), .ZN(n665) );
  NAND2_X4 U546 ( .A1(n2088), .A2(n1369), .ZN(n666) );
  XOR2_X2 U547 ( .A(n516), .B(n670), .Z(product[4]) );
  OAI21_X4 U548 ( .B1(n670), .B2(n668), .A(n669), .ZN(n667) );
  NAND2_X4 U549 ( .A1(n713), .A2(n669), .ZN(n516) );
  NOR2_X4 U551 ( .A1(n1371), .A2(n2089), .ZN(n668) );
  NAND2_X4 U552 ( .A1(n1371), .A2(n2089), .ZN(n669) );
  XNOR2_X2 U553 ( .A(n517), .B(n675), .ZN(product[3]) );
  AOI21_X4 U554 ( .B1(n675), .B2(n714), .A(n672), .ZN(n670) );
  NAND2_X4 U557 ( .A1(n714), .A2(n674), .ZN(n517) );
  XOR2_X2 U561 ( .A(n676), .B(n677), .Z(product[2]) );
  NOR2_X4 U562 ( .A1(n676), .A2(n677), .ZN(n675) );
  XNOR2_X2 U564 ( .A(n679), .B(n680), .ZN(product[1]) );
  NAND2_X4 U565 ( .A1(n678), .A2(n680), .ZN(n677) );
  FA_X1 U576 ( .A(n1721), .B(n1745), .CI(n723), .CO(n719), .S(n720) );
  FA_X1 U577 ( .A(n727), .B(n1722), .CI(n1746), .CO(n721), .S(n722) );
  FA_X1 U579 ( .A(n1747), .B(n727), .CI(n730), .CO(n725), .S(n726) );
  FA_X1 U581 ( .A(n734), .B(n1748), .CI(n731), .CO(n728), .S(n729) );
  FA_X1 U582 ( .A(n736), .B(n1779), .CI(n1723), .CO(n730), .S(n731) );
  FA_X1 U583 ( .A(n740), .B(n1749), .CI(n735), .CO(n732), .S(n733) );
  FA_X1 U584 ( .A(n742), .B(n1724), .CI(n1780), .CO(n734), .S(n735) );
  FA_X1 U586 ( .A(n741), .B(n747), .CI(n745), .CO(n738), .S(n739) );
  FA_X1 U587 ( .A(n1781), .B(n742), .CI(n1750), .CO(n740), .S(n741) );
  FA_X1 U589 ( .A(n751), .B(n748), .CI(n746), .CO(n743), .S(n744) );
  FA_X1 U590 ( .A(n1751), .B(n1782), .CI(n753), .CO(n745), .S(n746) );
  FA_X1 U591 ( .A(n755), .B(n1814), .CI(n1725), .CO(n747), .S(n748) );
  FA_X1 U592 ( .A(n759), .B(n754), .CI(n752), .CO(n749), .S(n750) );
  FA_X1 U593 ( .A(n1752), .B(n1783), .CI(n761), .CO(n751), .S(n752) );
  FA_X1 U594 ( .A(n763), .B(n1726), .CI(n1815), .CO(n753), .S(n754) );
  FA_X1 U596 ( .A(n766), .B(n762), .CI(n760), .CO(n757), .S(n758) );
  FA_X1 U597 ( .A(n770), .B(n1753), .CI(n768), .CO(n759), .S(n760) );
  FA_X1 U598 ( .A(n1816), .B(n763), .CI(n1784), .CO(n761), .S(n762) );
  FA_X1 U600 ( .A(n774), .B(n769), .CI(n767), .CO(n764), .S(n765) );
  FA_X1 U601 ( .A(n771), .B(n778), .CI(n776), .CO(n766), .S(n767) );
  FA_X1 U602 ( .A(n1785), .B(n1754), .CI(n1817), .CO(n768), .S(n769) );
  FA_X1 U603 ( .A(n780), .B(n1849), .CI(n1727), .CO(n770), .S(n771) );
  FA_X1 U604 ( .A(n784), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U605 ( .A(n779), .B(n788), .CI(n786), .CO(n774), .S(n775) );
  FA_X1 U606 ( .A(n1786), .B(n1755), .CI(n1818), .CO(n776), .S(n777) );
  FA_X1 U607 ( .A(n790), .B(n1728), .CI(n1850), .CO(n778), .S(n779) );
  FA_X1 U609 ( .A(n793), .B(n787), .CI(n785), .CO(n782), .S(n783) );
  FA_X1 U610 ( .A(n789), .B(n797), .CI(n795), .CO(n784), .S(n785) );
  FA_X1 U611 ( .A(n1787), .B(n1819), .CI(n799), .CO(n786), .S(n787) );
  FA_X1 U612 ( .A(n1851), .B(n790), .CI(n1756), .CO(n788), .S(n789) );
  FA_X1 U614 ( .A(n803), .B(n796), .CI(n794), .CO(n791), .S(n792) );
  FA_X1 U615 ( .A(n798), .B(n807), .CI(n805), .CO(n793), .S(n794) );
  FA_X1 U616 ( .A(n809), .B(n1820), .CI(n800), .CO(n795), .S(n796) );
  FA_X1 U617 ( .A(n1852), .B(n1757), .CI(n1788), .CO(n797), .S(n798) );
  FA_X1 U618 ( .A(n811), .B(n1884), .CI(n1729), .CO(n799), .S(n800) );
  FA_X1 U619 ( .A(n815), .B(n806), .CI(n804), .CO(n801), .S(n802) );
  FA_X1 U620 ( .A(n808), .B(n819), .CI(n817), .CO(n803), .S(n804) );
  FA_X1 U621 ( .A(n821), .B(n1758), .CI(n810), .CO(n805), .S(n806) );
  FA_X1 U622 ( .A(n1853), .B(n1789), .CI(n1821), .CO(n807), .S(n808) );
  FA_X1 U623 ( .A(n823), .B(n1730), .CI(n1885), .CO(n809), .S(n810) );
  FA_X1 U625 ( .A(n826), .B(n818), .CI(n816), .CO(n813), .S(n814) );
  FA_X1 U626 ( .A(n820), .B(n822), .CI(n828), .CO(n815), .S(n816) );
  FA_X1 U627 ( .A(n832), .B(n1759), .CI(n830), .CO(n817), .S(n818) );
  FA_X1 U628 ( .A(n1822), .B(n1790), .CI(n1854), .CO(n819), .S(n820) );
  FA_X1 U629 ( .A(n834), .B(n823), .CI(n1886), .CO(n821), .S(n822) );
  FA_X1 U631 ( .A(n838), .B(n829), .CI(n827), .CO(n824), .S(n825) );
  FA_X1 U632 ( .A(n842), .B(n833), .CI(n840), .CO(n826), .S(n827) );
  FA_X1 U633 ( .A(n844), .B(n846), .CI(n831), .CO(n828), .S(n829) );
  FA_X1 U634 ( .A(n1823), .B(n1760), .CI(n1887), .CO(n830), .S(n831) );
  FA_X1 U635 ( .A(n1855), .B(n1791), .CI(n835), .CO(n832), .S(n833) );
  FA_X1 U636 ( .A(n848), .B(n1919), .CI(n1731), .CO(n834), .S(n835) );
  FA_X1 U637 ( .A(n852), .B(n841), .CI(n839), .CO(n836), .S(n837) );
  FA_X1 U638 ( .A(n843), .B(n856), .CI(n854), .CO(n838), .S(n839) );
  FA_X1 U639 ( .A(n858), .B(n847), .CI(n845), .CO(n840), .S(n841) );
  FA_X1 U640 ( .A(n1761), .B(n1824), .CI(n860), .CO(n842), .S(n843) );
  FA_X1 U641 ( .A(n1888), .B(n1792), .CI(n1856), .CO(n844), .S(n845) );
  FA_X1 U642 ( .A(n1732), .B(n862), .CI(n1920), .CO(n846), .S(n847) );
  FA_X1 U644 ( .A(n865), .B(n855), .CI(n853), .CO(n850), .S(n851) );
  FA_X1 U645 ( .A(n857), .B(n869), .CI(n867), .CO(n852), .S(n853) );
  FA_X1 U646 ( .A(n861), .B(n871), .CI(n859), .CO(n854), .S(n855) );
  FA_X1 U647 ( .A(n1857), .B(n1762), .CI(n873), .CO(n856), .S(n857) );
  FA_X1 U648 ( .A(n1889), .B(n1793), .CI(n875), .CO(n858), .S(n859) );
  FA_X1 U649 ( .A(n1921), .B(n862), .CI(n1825), .CO(n860), .S(n861) );
  FA_X1 U651 ( .A(n879), .B(n868), .CI(n866), .CO(n863), .S(n864) );
  FA_X1 U652 ( .A(n870), .B(n883), .CI(n881), .CO(n865), .S(n866) );
  FA_X1 U653 ( .A(n874), .B(n885), .CI(n872), .CO(n867), .S(n868) );
  FA_X1 U654 ( .A(n889), .B(n876), .CI(n887), .CO(n869), .S(n870) );
  FA_X1 U655 ( .A(n1858), .B(n1922), .CI(n1890), .CO(n871), .S(n872) );
  FA_X1 U656 ( .A(n1826), .B(n1763), .CI(n1794), .CO(n873), .S(n874) );
  FA_X1 U657 ( .A(n891), .B(n1954), .CI(n1733), .CO(n875), .S(n876) );
  FA_X1 U658 ( .A(n895), .B(n882), .CI(n880), .CO(n877), .S(n878) );
  FA_X1 U659 ( .A(n884), .B(n899), .CI(n897), .CO(n879), .S(n880) );
  FA_X1 U660 ( .A(n888), .B(n901), .CI(n886), .CO(n881), .S(n882) );
  FA_X1 U661 ( .A(n890), .B(n905), .CI(n903), .CO(n883), .S(n884) );
  FA_X1 U662 ( .A(n1891), .B(n1859), .CI(n1923), .CO(n885), .S(n886) );
  FA_X1 U663 ( .A(n1827), .B(n1764), .CI(n1795), .CO(n887), .S(n888) );
  FA_X1 U664 ( .A(n907), .B(n892), .CI(n1955), .CO(n889), .S(n890) );
  FA_X1 U666 ( .A(n911), .B(n898), .CI(n896), .CO(n893), .S(n894) );
  FA_X1 U667 ( .A(n900), .B(n915), .CI(n913), .CO(n895), .S(n896) );
  FA_X1 U668 ( .A(n904), .B(n917), .CI(n902), .CO(n897), .S(n898) );
  FA_X1 U669 ( .A(n921), .B(n906), .CI(n919), .CO(n899), .S(n900) );
  FA_X1 U670 ( .A(n1892), .B(n1796), .CI(n1924), .CO(n901), .S(n902) );
  FA_X1 U671 ( .A(n1828), .B(n1956), .CI(n1860), .CO(n903), .S(n904) );
  FA_X1 U672 ( .A(n908), .B(n1734), .CI(n923), .CO(n905), .S(n906) );
  FA_X1 U674 ( .A(n927), .B(n914), .CI(n912), .CO(n909), .S(n910) );
  FA_X1 U675 ( .A(n916), .B(n931), .CI(n929), .CO(n911), .S(n912) );
  FA_X1 U676 ( .A(n920), .B(n933), .CI(n918), .CO(n913), .S(n914) );
  FA_X1 U677 ( .A(n935), .B(n937), .CI(n922), .CO(n915), .S(n916) );
  FA_X1 U678 ( .A(n1893), .B(n1829), .CI(n1957), .CO(n917), .S(n918) );
  FA_X1 U679 ( .A(n1925), .B(n1861), .CI(n939), .CO(n919), .S(n920) );
  FA_X1 U680 ( .A(n1765), .B(n1797), .CI(n924), .CO(n921), .S(n922) );
  FA_X1 U681 ( .A(n941), .B(n1989), .CI(n1735), .CO(n923), .S(n924) );
  FA_X1 U682 ( .A(n945), .B(n930), .CI(n928), .CO(n925), .S(n926) );
  FA_X1 U683 ( .A(n932), .B(n949), .CI(n947), .CO(n927), .S(n928) );
  FA_X1 U684 ( .A(n951), .B(n936), .CI(n934), .CO(n929), .S(n930) );
  FA_X1 U685 ( .A(n953), .B(n955), .CI(n938), .CO(n931), .S(n932) );
  FA_X1 U686 ( .A(n957), .B(n1894), .CI(n940), .CO(n933), .S(n934) );
  FA_X1 U687 ( .A(n1926), .B(n1830), .CI(n1958), .CO(n935), .S(n936) );
  FA_X1 U688 ( .A(n1798), .B(n1990), .CI(n1862), .CO(n937), .S(n938) );
  FA_X1 U689 ( .A(n1736), .B(n959), .CI(n1766), .CO(n939), .S(n940) );
  FA_X1 U691 ( .A(n962), .B(n948), .CI(n946), .CO(n943), .S(n944) );
  FA_X1 U692 ( .A(n950), .B(n966), .CI(n964), .CO(n945), .S(n946) );
  FA_X1 U693 ( .A(n968), .B(n954), .CI(n952), .CO(n947), .S(n948) );
  FA_X1 U694 ( .A(n970), .B(n972), .CI(n956), .CO(n949), .S(n950) );
  FA_X1 U695 ( .A(n974), .B(n1895), .CI(n958), .CO(n951), .S(n952) );
  FA_X1 U696 ( .A(n1927), .B(n1831), .CI(n1959), .CO(n953), .S(n954) );
  FA_X1 U697 ( .A(n1767), .B(n1991), .CI(n1863), .CO(n955), .S(n956) );
  FA_X1 U698 ( .A(n1799), .B(n959), .CI(n976), .CO(n957), .S(n958) );
  FA_X1 U700 ( .A(n980), .B(n965), .CI(n963), .CO(n960), .S(n961) );
  FA_X1 U701 ( .A(n967), .B(n969), .CI(n982), .CO(n962), .S(n963) );
  FA_X1 U702 ( .A(n986), .B(n971), .CI(n984), .CO(n964), .S(n965) );
  FA_X1 U703 ( .A(n975), .B(n988), .CI(n973), .CO(n966), .S(n967) );
  FA_X1 U704 ( .A(n992), .B(n1960), .CI(n990), .CO(n968), .S(n969) );
  FA_X1 U705 ( .A(n1928), .B(n1992), .CI(n994), .CO(n970), .S(n971) );
  FA_X1 U706 ( .A(n1896), .B(n977), .CI(n1864), .CO(n972), .S(n973) );
  FA_X1 U707 ( .A(n1832), .B(n1768), .CI(n1800), .CO(n974), .S(n975) );
  FA_X1 U708 ( .A(n2024), .B(n2059), .CI(n1737), .CO(n976), .S(n977) );
  FA_X1 U709 ( .A(n998), .B(n983), .CI(n981), .CO(n978), .S(n979) );
  FA_X1 U710 ( .A(n985), .B(n987), .CI(n1000), .CO(n980), .S(n981) );
  FA_X1 U711 ( .A(n1004), .B(n989), .CI(n1002), .CO(n982), .S(n983) );
  FA_X1 U712 ( .A(n993), .B(n1006), .CI(n991), .CO(n984), .S(n985) );
  FA_X1 U713 ( .A(n1010), .B(n995), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U714 ( .A(n1865), .B(n1929), .CI(n1961), .CO(n988), .S(n989) );
  FA_X1 U715 ( .A(n1897), .B(n1012), .CI(n1993), .CO(n990), .S(n991) );
  FA_X1 U716 ( .A(n2025), .B(n1769), .CI(n1833), .CO(n992), .S(n993) );
  FA_X1 U717 ( .A(n1738), .B(n262), .CI(n1801), .CO(n994), .S(n995) );
  FA_X1 U718 ( .A(n1016), .B(n1001), .CI(n999), .CO(n996), .S(n997) );
  FA_X1 U719 ( .A(n1003), .B(n1005), .CI(n1018), .CO(n998), .S(n999) );
  FA_X1 U720 ( .A(n1022), .B(n1009), .CI(n1020), .CO(n1000), .S(n1001) );
  FA_X1 U721 ( .A(n1011), .B(n1024), .CI(n1007), .CO(n1002), .S(n1003) );
  FA_X1 U722 ( .A(n1028), .B(n1013), .CI(n1026), .CO(n1004), .S(n1005) );
  FA_X1 U723 ( .A(n1866), .B(n1930), .CI(n1962), .CO(n1006), .S(n1007) );
  FA_X1 U724 ( .A(n1994), .B(n1898), .CI(n1030), .CO(n1008), .S(n1009) );
  FA_X1 U725 ( .A(n2026), .B(n1834), .CI(n1802), .CO(n1010), .S(n1011) );
  FA_X1 U726 ( .A(n1739), .B(n262), .CI(n1770), .CO(n1012), .S(n1013) );
  FA_X1 U727 ( .A(n1034), .B(n1019), .CI(n1017), .CO(n1014), .S(n1015) );
  FA_X1 U728 ( .A(n1021), .B(n1023), .CI(n1036), .CO(n1016), .S(n1017) );
  FA_X1 U729 ( .A(n1040), .B(n1027), .CI(n1038), .CO(n1018), .S(n1019) );
  FA_X1 U730 ( .A(n1029), .B(n1042), .CI(n1025), .CO(n1020), .S(n1021) );
  FA_X1 U731 ( .A(n1046), .B(n1031), .CI(n1044), .CO(n1022), .S(n1023) );
  FA_X1 U732 ( .A(n1963), .B(n1899), .CI(n1995), .CO(n1024), .S(n1025) );
  FA_X1 U733 ( .A(n2027), .B(n1931), .CI(n1048), .CO(n1026), .S(n1027) );
  FA_X1 U734 ( .A(n1867), .B(n1803), .CI(n1835), .CO(n1028), .S(n1029) );
  FA_X1 U735 ( .A(n1740), .B(n262), .CI(n1771), .CO(n1030), .S(n1031) );
  FA_X1 U736 ( .A(n1052), .B(n1037), .CI(n1035), .CO(n1032), .S(n1033) );
  FA_X1 U737 ( .A(n1039), .B(n1041), .CI(n1054), .CO(n1034), .S(n1035) );
  FA_X1 U738 ( .A(n1058), .B(n1045), .CI(n1056), .CO(n1036), .S(n1037) );
  FA_X1 U739 ( .A(n1047), .B(n1060), .CI(n1043), .CO(n1038), .S(n1039) );
  FA_X1 U740 ( .A(n1064), .B(n1049), .CI(n1062), .CO(n1040), .S(n1041) );
  FA_X1 U741 ( .A(n1900), .B(n1964), .CI(n1066), .CO(n1042), .S(n1043) );
  FA_X1 U742 ( .A(n2028), .B(n1932), .CI(n1996), .CO(n1044), .S(n1045) );
  FA_X1 U743 ( .A(n2060), .B(n1836), .CI(n1868), .CO(n1046), .S(n1047) );
  FA_X1 U744 ( .A(n1772), .B(n1741), .CI(n1804), .CO(n1048), .S(n1049) );
  FA_X1 U745 ( .A(n1070), .B(n1055), .CI(n1053), .CO(n1050), .S(n1051) );
  FA_X1 U746 ( .A(n1057), .B(n1059), .CI(n1072), .CO(n1052), .S(n1053) );
  FA_X1 U747 ( .A(n1076), .B(n1063), .CI(n1074), .CO(n1054), .S(n1055) );
  FA_X1 U748 ( .A(n1065), .B(n1078), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U749 ( .A(n1067), .B(n1082), .CI(n1080), .CO(n1058), .S(n1059) );
  FA_X1 U750 ( .A(n1933), .B(n1965), .CI(n1997), .CO(n1060), .S(n1061) );
  FA_X1 U751 ( .A(n2029), .B(n1901), .CI(n1084), .CO(n1062), .S(n1063) );
  FA_X1 U752 ( .A(n2061), .B(n1869), .CI(n1837), .CO(n1064), .S(n1065) );
  FA_X1 U753 ( .A(n1773), .B(n1742), .CI(n1805), .CO(n1066), .S(n1067) );
  FA_X1 U754 ( .A(n1088), .B(n1073), .CI(n1071), .CO(n1068), .S(n1069) );
  FA_X1 U755 ( .A(n1075), .B(n1092), .CI(n1090), .CO(n1070), .S(n1071) );
  FA_X1 U756 ( .A(n1079), .B(n1094), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U757 ( .A(n1096), .B(n1098), .CI(n1081), .CO(n1074), .S(n1075) );
  FA_X1 U758 ( .A(n1085), .B(n1100), .CI(n1083), .CO(n1076), .S(n1077) );
  FA_X1 U759 ( .A(n1998), .B(n2062), .CI(n2030), .CO(n1078), .S(n1079) );
  FA_X1 U760 ( .A(n1966), .B(n1870), .CI(n1934), .CO(n1080), .S(n1081) );
  FA_X1 U761 ( .A(n1102), .B(n1838), .CI(n1902), .CO(n1082), .S(n1083) );
  FA_X1 U762 ( .A(n1774), .B(n1743), .CI(n1806), .CO(n1084), .S(n1085) );
  FA_X1 U763 ( .A(n1106), .B(n1091), .CI(n1089), .CO(n1086), .S(n1087) );
  FA_X1 U764 ( .A(n1108), .B(n1110), .CI(n1093), .CO(n1088), .S(n1089) );
  FA_X1 U765 ( .A(n1097), .B(n1099), .CI(n1095), .CO(n1090), .S(n1091) );
  FA_X1 U766 ( .A(n1114), .B(n1116), .CI(n1112), .CO(n1092), .S(n1093) );
  FA_X1 U767 ( .A(n1118), .B(n1999), .CI(n1101), .CO(n1094), .S(n1095) );
  FA_X1 U768 ( .A(n2063), .B(n1935), .CI(n2031), .CO(n1096), .S(n1097) );
  FA_X1 U769 ( .A(n1903), .B(n1103), .CI(n1967), .CO(n1098), .S(n1099) );
  FA_X1 U770 ( .A(n1871), .B(n1807), .CI(n1839), .CO(n1100), .S(n1101) );
  FA_X1 U771 ( .A(n1775), .B(n1744), .CI(n1120), .CO(n1102), .S(n1103) );
  FA_X1 U772 ( .A(n1124), .B(n1109), .CI(n1107), .CO(n1104), .S(n1105) );
  FA_X1 U773 ( .A(n1126), .B(n1128), .CI(n1111), .CO(n1106), .S(n1107) );
  FA_X1 U774 ( .A(n1115), .B(n1117), .CI(n1113), .CO(n1108), .S(n1109) );
  FA_X1 U775 ( .A(n1132), .B(n1119), .CI(n1130), .CO(n1110), .S(n1111) );
  FA_X1 U776 ( .A(n2064), .B(n2000), .CI(n1134), .CO(n1112), .S(n1113) );
  FA_X1 U777 ( .A(n2032), .B(n1936), .CI(n1136), .CO(n1114), .S(n1115) );
  FA_X1 U778 ( .A(n1872), .B(n1904), .CI(n1968), .CO(n1116), .S(n1117) );
  FA_X1 U779 ( .A(n1808), .B(n1121), .CI(n1840), .CO(n1118), .S(n1119) );
  HA_X1 U780 ( .A(n1776), .B(n1138), .CO(n1120), .S(n1121) );
  FA_X1 U781 ( .A(n1142), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U782 ( .A(n1129), .B(n1146), .CI(n1144), .CO(n1124), .S(n1125) );
  FA_X1 U783 ( .A(n1133), .B(n1148), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U784 ( .A(n1135), .B(n1137), .CI(n1150), .CO(n1128), .S(n1129) );
  FA_X1 U785 ( .A(n2033), .B(n2065), .CI(n1152), .CO(n1130), .S(n1131) );
  FA_X1 U786 ( .A(n2001), .B(n1905), .CI(n1969), .CO(n1132), .S(n1133) );
  FA_X1 U787 ( .A(n1154), .B(n1873), .CI(n1937), .CO(n1134), .S(n1135) );
  FA_X1 U788 ( .A(n1139), .B(n1809), .CI(n1841), .CO(n1136), .S(n1137) );
  HA_X1 U789 ( .A(n1156), .B(n1777), .CO(n1138), .S(n1139) );
  FA_X1 U790 ( .A(n1160), .B(n1145), .CI(n1143), .CO(n1140), .S(n1141) );
  FA_X1 U791 ( .A(n1147), .B(n1149), .CI(n1162), .CO(n1142), .S(n1143) );
  FA_X1 U792 ( .A(n1164), .B(n1166), .CI(n1151), .CO(n1144), .S(n1145) );
  FA_X1 U793 ( .A(n1153), .B(n2002), .CI(n1168), .CO(n1146), .S(n1147) );
  FA_X1 U794 ( .A(n1170), .B(n2034), .CI(n2066), .CO(n1148), .S(n1149) );
  FA_X1 U795 ( .A(n1938), .B(n1155), .CI(n1970), .CO(n1150), .S(n1151) );
  FA_X1 U796 ( .A(n1874), .B(n1842), .CI(n1906), .CO(n1152), .S(n1153) );
  FA_X1 U797 ( .A(n1810), .B(n1157), .CI(n1172), .CO(n1154), .S(n1155) );
  HA_X1 U798 ( .A(n289), .B(n1778), .CO(n1156), .S(n1157) );
  FA_X1 U799 ( .A(n1176), .B(n1163), .CI(n1161), .CO(n1158), .S(n1159) );
  FA_X1 U800 ( .A(n1165), .B(n1167), .CI(n1178), .CO(n1160), .S(n1161) );
  FA_X1 U801 ( .A(n1169), .B(n1182), .CI(n1180), .CO(n1162), .S(n1163) );
  FA_X1 U802 ( .A(n1184), .B(n2003), .CI(n1171), .CO(n1164), .S(n1165) );
  FA_X1 U803 ( .A(n2067), .B(n2035), .CI(n1186), .CO(n1166), .S(n1167) );
  FA_X1 U804 ( .A(n1907), .B(n1939), .CI(n1971), .CO(n1168), .S(n1169) );
  FA_X1 U805 ( .A(n1843), .B(n1173), .CI(n1875), .CO(n1170), .S(n1171) );
  HA_X1 U806 ( .A(n1811), .B(n1188), .CO(n1172), .S(n1173) );
  FA_X1 U807 ( .A(n1192), .B(n1179), .CI(n1177), .CO(n1174), .S(n1175) );
  FA_X1 U808 ( .A(n1181), .B(n1183), .CI(n1194), .CO(n1176), .S(n1177) );
  FA_X1 U809 ( .A(n1198), .B(n1185), .CI(n1196), .CO(n1178), .S(n1179) );
  FA_X1 U810 ( .A(n1200), .B(n2068), .CI(n1187), .CO(n1180), .S(n1181) );
  FA_X1 U811 ( .A(n2004), .B(n1940), .CI(n2036), .CO(n1182), .S(n1183) );
  FA_X1 U812 ( .A(n1202), .B(n1908), .CI(n1972), .CO(n1184), .S(n1185) );
  FA_X1 U813 ( .A(n1189), .B(n1844), .CI(n1876), .CO(n1186), .S(n1187) );
  HA_X1 U814 ( .A(n1204), .B(n1812), .CO(n1188), .S(n1189) );
  FA_X1 U815 ( .A(n1208), .B(n1195), .CI(n1193), .CO(n1190), .S(n1191) );
  FA_X1 U816 ( .A(n1197), .B(n1199), .CI(n1210), .CO(n1192), .S(n1193) );
  FA_X1 U817 ( .A(n1214), .B(n1201), .CI(n1212), .CO(n1194), .S(n1195) );
  FA_X1 U818 ( .A(n2037), .B(n2069), .CI(n1216), .CO(n1196), .S(n1197) );
  FA_X1 U819 ( .A(n1973), .B(n1203), .CI(n2005), .CO(n1198), .S(n1199) );
  FA_X1 U820 ( .A(n1941), .B(n1877), .CI(n1909), .CO(n1200), .S(n1201) );
  FA_X1 U821 ( .A(n1845), .B(n1205), .CI(n1218), .CO(n1202), .S(n1203) );
  HA_X1 U822 ( .A(n286), .B(n1813), .CO(n1204), .S(n1205) );
  FA_X1 U823 ( .A(n1222), .B(n1211), .CI(n1209), .CO(n1206), .S(n1207) );
  FA_X1 U824 ( .A(n1213), .B(n1215), .CI(n1224), .CO(n1208), .S(n1209) );
  FA_X1 U825 ( .A(n1217), .B(n1228), .CI(n1226), .CO(n1210), .S(n1211) );
  FA_X1 U826 ( .A(n2038), .B(n2070), .CI(n1230), .CO(n1212), .S(n1213) );
  FA_X1 U827 ( .A(n1942), .B(n1974), .CI(n2006), .CO(n1214), .S(n1215) );
  FA_X1 U828 ( .A(n1878), .B(n1219), .CI(n1910), .CO(n1216), .S(n1217) );
  HA_X1 U829 ( .A(n1846), .B(n1232), .CO(n1218), .S(n1219) );
  FA_X1 U830 ( .A(n1236), .B(n1225), .CI(n1223), .CO(n1220), .S(n1221) );
  FA_X1 U831 ( .A(n1227), .B(n1240), .CI(n1238), .CO(n1222), .S(n1223) );
  FA_X1 U832 ( .A(n1231), .B(n1242), .CI(n1229), .CO(n1224), .S(n1225) );
  FA_X1 U833 ( .A(n2071), .B(n1975), .CI(n2039), .CO(n1226), .S(n1227) );
  FA_X1 U834 ( .A(n1244), .B(n1943), .CI(n2007), .CO(n1228), .S(n1229) );
  FA_X1 U835 ( .A(n1233), .B(n1879), .CI(n1911), .CO(n1230), .S(n1231) );
  HA_X1 U836 ( .A(n1246), .B(n1847), .CO(n1232), .S(n1233) );
  FA_X1 U837 ( .A(n1250), .B(n1239), .CI(n1237), .CO(n1234), .S(n1235) );
  FA_X1 U838 ( .A(n1252), .B(n1254), .CI(n1241), .CO(n1236), .S(n1237) );
  FA_X1 U839 ( .A(n1256), .B(n2040), .CI(n1243), .CO(n1238), .S(n1239) );
  FA_X1 U840 ( .A(n2008), .B(n1245), .CI(n2072), .CO(n1240), .S(n1241) );
  FA_X1 U841 ( .A(n1944), .B(n1912), .CI(n1976), .CO(n1242), .S(n1243) );
  FA_X1 U842 ( .A(n1880), .B(n1247), .CI(n1258), .CO(n1244), .S(n1245) );
  HA_X1 U843 ( .A(n283), .B(n1848), .CO(n1246), .S(n1247) );
  FA_X1 U844 ( .A(n1262), .B(n1253), .CI(n1251), .CO(n1248), .S(n1249) );
  FA_X1 U845 ( .A(n1264), .B(n1257), .CI(n1255), .CO(n1250), .S(n1251) );
  FA_X1 U846 ( .A(n1268), .B(n2041), .CI(n1266), .CO(n1252), .S(n1253) );
  FA_X1 U847 ( .A(n1977), .B(n2009), .CI(n2073), .CO(n1254), .S(n1255) );
  FA_X1 U848 ( .A(n1913), .B(n1259), .CI(n1945), .CO(n1256), .S(n1257) );
  HA_X1 U849 ( .A(n1881), .B(n1270), .CO(n1258), .S(n1259) );
  FA_X1 U850 ( .A(n1274), .B(n1265), .CI(n1263), .CO(n1260), .S(n1261) );
  FA_X1 U851 ( .A(n1267), .B(n1269), .CI(n1276), .CO(n1262), .S(n1263) );
  FA_X1 U852 ( .A(n2074), .B(n2010), .CI(n1278), .CO(n1264), .S(n1265) );
  FA_X1 U853 ( .A(n1280), .B(n1978), .CI(n2042), .CO(n1266), .S(n1267) );
  FA_X1 U854 ( .A(n1271), .B(n1914), .CI(n1946), .CO(n1268), .S(n1269) );
  HA_X1 U855 ( .A(n1282), .B(n1882), .CO(n1270), .S(n1271) );
  FA_X1 U856 ( .A(n1277), .B(n1286), .CI(n1275), .CO(n1272), .S(n1273) );
  FA_X1 U857 ( .A(n1279), .B(n1290), .CI(n1288), .CO(n1274), .S(n1275) );
  FA_X1 U858 ( .A(n2043), .B(n1281), .CI(n2075), .CO(n1276), .S(n1277) );
  FA_X1 U859 ( .A(n2011), .B(n1947), .CI(n1979), .CO(n1278), .S(n1279) );
  FA_X1 U860 ( .A(n1915), .B(n1283), .CI(n1292), .CO(n1280), .S(n1281) );
  HA_X1 U861 ( .A(n280), .B(n1883), .CO(n1282), .S(n1283) );
  FA_X1 U862 ( .A(n1296), .B(n1289), .CI(n1287), .CO(n1284), .S(n1285) );
  FA_X1 U863 ( .A(n1298), .B(n1300), .CI(n1291), .CO(n1286), .S(n1287) );
  FA_X1 U864 ( .A(n2012), .B(n2044), .CI(n2076), .CO(n1288), .S(n1289) );
  FA_X1 U865 ( .A(n1948), .B(n1293), .CI(n1980), .CO(n1290), .S(n1291) );
  HA_X1 U866 ( .A(n1916), .B(n1302), .CO(n1292), .S(n1293) );
  FA_X1 U867 ( .A(n1306), .B(n1299), .CI(n1297), .CO(n1294), .S(n1295) );
  FA_X1 U868 ( .A(n1308), .B(n2045), .CI(n1301), .CO(n1296), .S(n1297) );
  FA_X1 U869 ( .A(n1310), .B(n2013), .CI(n2077), .CO(n1298), .S(n1299) );
  FA_X1 U870 ( .A(n1303), .B(n1949), .CI(n1981), .CO(n1300), .S(n1301) );
  HA_X1 U871 ( .A(n1312), .B(n1917), .CO(n1302), .S(n1303) );
  FA_X1 U872 ( .A(n1316), .B(n1309), .CI(n1307), .CO(n1304), .S(n1305) );
  FA_X1 U873 ( .A(n2078), .B(n1311), .CI(n1318), .CO(n1306), .S(n1307) );
  FA_X1 U874 ( .A(n2046), .B(n1982), .CI(n2014), .CO(n1308), .S(n1309) );
  FA_X1 U875 ( .A(n1950), .B(n1313), .CI(n1320), .CO(n1310), .S(n1311) );
  HA_X1 U876 ( .A(n277), .B(n1918), .CO(n1312), .S(n1313) );
  FA_X1 U877 ( .A(n1324), .B(n1319), .CI(n1317), .CO(n1314), .S(n1315) );
  FA_X1 U878 ( .A(n2047), .B(n2079), .CI(n1326), .CO(n1316), .S(n1317) );
  FA_X1 U879 ( .A(n1983), .B(n1321), .CI(n2015), .CO(n1318), .S(n1319) );
  HA_X1 U880 ( .A(n1951), .B(n1328), .CO(n1320), .S(n1321) );
  FA_X1 U881 ( .A(n1327), .B(n1332), .CI(n1325), .CO(n1322), .S(n1323) );
  FA_X1 U882 ( .A(n1334), .B(n2048), .CI(n2080), .CO(n1324), .S(n1325) );
  FA_X1 U883 ( .A(n1329), .B(n1984), .CI(n2016), .CO(n1326), .S(n1327) );
  HA_X1 U884 ( .A(n1336), .B(n1952), .CO(n1328), .S(n1329) );
  FA_X1 U885 ( .A(n1340), .B(n1335), .CI(n1333), .CO(n1330), .S(n1331) );
  FA_X1 U886 ( .A(n2081), .B(n2017), .CI(n2049), .CO(n1332), .S(n1333) );
  FA_X1 U887 ( .A(n1985), .B(n1337), .CI(n1342), .CO(n1334), .S(n1335) );
  HA_X1 U888 ( .A(n274), .B(n1953), .CO(n1336), .S(n1337) );
  FA_X1 U889 ( .A(n1346), .B(n2082), .CI(n1341), .CO(n1338), .S(n1339) );
  FA_X1 U890 ( .A(n2018), .B(n1343), .CI(n2050), .CO(n1340), .S(n1341) );
  HA_X1 U891 ( .A(n1986), .B(n1348), .CO(n1342), .S(n1343) );
  FA_X1 U892 ( .A(n1352), .B(n2083), .CI(n1347), .CO(n1344), .S(n1345) );
  FA_X1 U893 ( .A(n1349), .B(n2019), .CI(n2051), .CO(n1346), .S(n1347) );
  HA_X1 U894 ( .A(n1354), .B(n1987), .CO(n1348), .S(n1349) );
  FA_X1 U895 ( .A(n2084), .B(n2052), .CI(n1353), .CO(n1350), .S(n1351) );
  FA_X1 U896 ( .A(n2020), .B(n1355), .CI(n1358), .CO(n1352), .S(n1353) );
  HA_X1 U897 ( .A(n271), .B(n1988), .CO(n1354), .S(n1355) );
  FA_X1 U898 ( .A(n2053), .B(n1359), .CI(n2085), .CO(n1356), .S(n1357) );
  HA_X1 U899 ( .A(n2021), .B(n1362), .CO(n1358), .S(n1359) );
  FA_X1 U900 ( .A(n1363), .B(n2054), .CI(n2086), .CO(n1360), .S(n1361) );
  HA_X1 U901 ( .A(n1366), .B(n2022), .CO(n1362), .S(n1363) );
  FA_X1 U902 ( .A(n2055), .B(n1367), .CI(n1368), .CO(n1364), .S(n1365) );
  HA_X1 U903 ( .A(n268), .B(n2023), .CO(n1366), .S(n1367) );
  HA_X1 U904 ( .A(n2056), .B(n1370), .CO(n1368), .S(n1369) );
  HA_X1 U905 ( .A(n1372), .B(n2057), .CO(n1370), .S(n1371) );
  HA_X1 U906 ( .A(n265), .B(n2058), .CO(n1372), .S(n1373) );
  OAI21_X4 U907 ( .B1(n2808), .B2(n3161), .A(n2094), .ZN(n1720) );
  NAND2_X4 U908 ( .A1(n388), .A2(n484), .ZN(n2094) );
  OAI21_X4 U909 ( .B1(n2809), .B2(n3161), .A(n2095), .ZN(n717) );
  AOI21_X4 U910 ( .B1(n388), .B2(n481), .A(n1374), .ZN(n2095) );
  AND2_X4 U911 ( .A1(n333), .A2(n484), .ZN(n1374) );
  OAI21_X4 U912 ( .B1(n2810), .B2(n3161), .A(n2096), .ZN(n1721) );
  AOI222_X2 U913 ( .A1(n3131), .A2(n484), .B1(n333), .B2(n481), .C1(n388), 
        .C2(n478), .ZN(n2096) );
  OAI21_X4 U914 ( .B1(n2811), .B2(n3161), .A(n2097), .ZN(n1722) );
  AOI222_X2 U915 ( .A1(n3130), .A2(n481), .B1(n333), .B2(n478), .C1(n388), 
        .C2(n475), .ZN(n2097) );
  OAI21_X4 U916 ( .B1(n2812), .B2(n3161), .A(n2098), .ZN(n723) );
  AOI222_X2 U917 ( .A1(n3131), .A2(n478), .B1(n333), .B2(n475), .C1(n388), 
        .C2(n472), .ZN(n2098) );
  OAI21_X4 U918 ( .B1(n2813), .B2(n3161), .A(n2099), .ZN(n1723) );
  AOI222_X2 U919 ( .A1(n3130), .A2(n475), .B1(n333), .B2(n472), .C1(n388), 
        .C2(n469), .ZN(n2099) );
  OAI21_X4 U920 ( .B1(n2814), .B2(n3161), .A(n2100), .ZN(n1724) );
  AOI222_X2 U921 ( .A1(n3131), .A2(n472), .B1(n333), .B2(n469), .C1(n388), 
        .C2(n466), .ZN(n2100) );
  OAI21_X4 U922 ( .B1(n2815), .B2(n3161), .A(n2101), .ZN(n736) );
  AOI222_X2 U923 ( .A1(n3130), .A2(n469), .B1(n333), .B2(n466), .C1(n388), 
        .C2(n463), .ZN(n2101) );
  OAI21_X4 U924 ( .B1(n2816), .B2(n3161), .A(n2102), .ZN(n1725) );
  AOI222_X2 U925 ( .A1(n3131), .A2(n466), .B1(n333), .B2(n463), .C1(n388), 
        .C2(n460), .ZN(n2102) );
  OAI21_X4 U926 ( .B1(n2817), .B2(n3161), .A(n2103), .ZN(n1726) );
  AOI222_X2 U927 ( .A1(n3130), .A2(n463), .B1(n333), .B2(n460), .C1(n388), 
        .C2(n457), .ZN(n2103) );
  OAI21_X4 U928 ( .B1(n2818), .B2(n3161), .A(n2104), .ZN(n755) );
  AOI222_X2 U929 ( .A1(n3131), .A2(n460), .B1(n333), .B2(n457), .C1(n388), 
        .C2(n454), .ZN(n2104) );
  OAI21_X4 U930 ( .B1(n2819), .B2(n3161), .A(n2105), .ZN(n1727) );
  AOI222_X2 U931 ( .A1(n3130), .A2(n457), .B1(n333), .B2(n454), .C1(n388), 
        .C2(n451), .ZN(n2105) );
  OAI21_X4 U932 ( .B1(n2820), .B2(n3161), .A(n2106), .ZN(n1728) );
  AOI222_X2 U933 ( .A1(n3131), .A2(n454), .B1(n333), .B2(n451), .C1(n388), 
        .C2(n448), .ZN(n2106) );
  OAI21_X4 U934 ( .B1(n2821), .B2(n3161), .A(n2107), .ZN(n780) );
  AOI222_X2 U935 ( .A1(n3130), .A2(n451), .B1(n333), .B2(n448), .C1(n388), 
        .C2(n445), .ZN(n2107) );
  OAI21_X4 U936 ( .B1(n2822), .B2(n3161), .A(n2108), .ZN(n1729) );
  AOI222_X2 U937 ( .A1(n3131), .A2(n448), .B1(n333), .B2(n445), .C1(n388), 
        .C2(n442), .ZN(n2108) );
  OAI21_X4 U938 ( .B1(n2823), .B2(n3161), .A(n2109), .ZN(n1730) );
  AOI222_X2 U939 ( .A1(n3130), .A2(n445), .B1(n333), .B2(n442), .C1(n388), 
        .C2(n439), .ZN(n2109) );
  OAI21_X4 U940 ( .B1(n2824), .B2(n3161), .A(n2110), .ZN(n811) );
  AOI222_X2 U941 ( .A1(n3131), .A2(n442), .B1(n333), .B2(n439), .C1(n388), 
        .C2(n436), .ZN(n2110) );
  OAI21_X4 U942 ( .B1(n2825), .B2(n3161), .A(n2111), .ZN(n1731) );
  AOI222_X2 U943 ( .A1(n3130), .A2(n439), .B1(n333), .B2(n436), .C1(n388), 
        .C2(n433), .ZN(n2111) );
  OAI21_X4 U944 ( .B1(n2826), .B2(n3161), .A(n2112), .ZN(n1732) );
  AOI222_X2 U945 ( .A1(n3131), .A2(n436), .B1(n333), .B2(n433), .C1(n388), 
        .C2(n430), .ZN(n2112) );
  OAI21_X4 U946 ( .B1(n2827), .B2(n3161), .A(n2113), .ZN(n848) );
  AOI222_X2 U947 ( .A1(n3130), .A2(n433), .B1(n333), .B2(n430), .C1(n388), 
        .C2(n427), .ZN(n2113) );
  OAI21_X4 U948 ( .B1(n2828), .B2(n3161), .A(n2114), .ZN(n1733) );
  AOI222_X2 U949 ( .A1(n3131), .A2(n430), .B1(n333), .B2(n427), .C1(n388), 
        .C2(n424), .ZN(n2114) );
  OAI21_X4 U950 ( .B1(n2829), .B2(n3161), .A(n2115), .ZN(n891) );
  AOI222_X2 U951 ( .A1(n3130), .A2(n427), .B1(n333), .B2(n424), .C1(n388), 
        .C2(n421), .ZN(n2115) );
  OAI21_X4 U952 ( .B1(n2830), .B2(n3161), .A(n2116), .ZN(n1734) );
  AOI222_X2 U953 ( .A1(n3131), .A2(n424), .B1(n333), .B2(n421), .C1(n388), 
        .C2(n418), .ZN(n2116) );
  OAI21_X4 U954 ( .B1(n2831), .B2(n3161), .A(n2117), .ZN(n1735) );
  AOI222_X2 U955 ( .A1(n3131), .A2(n421), .B1(n333), .B2(n418), .C1(n388), 
        .C2(n415), .ZN(n2117) );
  OAI21_X4 U956 ( .B1(n2832), .B2(n3161), .A(n2118), .ZN(n1736) );
  AOI222_X2 U957 ( .A1(n3130), .A2(n418), .B1(n333), .B2(n415), .C1(n388), 
        .C2(n412), .ZN(n2118) );
  OAI21_X4 U958 ( .B1(n2833), .B2(n3161), .A(n2119), .ZN(n941) );
  AOI222_X2 U959 ( .A1(n3130), .A2(n415), .B1(n333), .B2(n412), .C1(n388), 
        .C2(n409), .ZN(n2119) );
  OAI21_X4 U960 ( .B1(n2834), .B2(n3160), .A(n2120), .ZN(n1737) );
  AOI222_X2 U961 ( .A1(n3130), .A2(n412), .B1(n333), .B2(n409), .C1(n388), 
        .C2(n406), .ZN(n2120) );
  OAI21_X4 U962 ( .B1(n2835), .B2(n3160), .A(n2121), .ZN(n1738) );
  AOI222_X2 U963 ( .A1(n3131), .A2(n409), .B1(n333), .B2(n406), .C1(n388), 
        .C2(n403), .ZN(n2121) );
  OAI21_X4 U964 ( .B1(n2836), .B2(n3160), .A(n2122), .ZN(n1739) );
  AOI222_X2 U965 ( .A1(n3131), .A2(n406), .B1(n333), .B2(n403), .C1(n388), 
        .C2(n400), .ZN(n2122) );
  OAI21_X4 U966 ( .B1(n2837), .B2(n3160), .A(n2123), .ZN(n1740) );
  AOI222_X2 U967 ( .A1(n3130), .A2(n403), .B1(n333), .B2(n400), .C1(n388), 
        .C2(n397), .ZN(n2123) );
  OAI21_X4 U968 ( .B1(n2838), .B2(n3160), .A(n2124), .ZN(n1741) );
  AOI222_X2 U969 ( .A1(n3131), .A2(n400), .B1(n333), .B2(n397), .C1(n388), 
        .C2(n393), .ZN(n2124) );
  OAI21_X4 U970 ( .B1(n2839), .B2(n3160), .A(n2125), .ZN(n1742) );
  AOI222_X2 U971 ( .A1(n3131), .A2(n397), .B1(n333), .B2(n393), .C1(n388), 
        .C2(n390), .ZN(n2125) );
  OAI21_X4 U972 ( .B1(n2840), .B2(n3160), .A(n2126), .ZN(n1743) );
  OAI21_X4 U974 ( .B1(n2841), .B2(n3160), .A(n2127), .ZN(n1744) );
  AND2_X4 U976 ( .A1(n3130), .A2(n390), .ZN(n1376) );
  XOR2_X2 U978 ( .A(n2128), .B(n289), .Z(n1746) );
  OAI21_X4 U979 ( .B1(n2808), .B2(n3158), .A(n2162), .ZN(n2128) );
  NAND2_X4 U980 ( .A1(n386), .A2(n484), .ZN(n2162) );
  XOR2_X2 U981 ( .A(n2129), .B(n289), .Z(n1747) );
  OAI21_X4 U982 ( .B1(n2809), .B2(n3158), .A(n2163), .ZN(n2129) );
  AOI21_X4 U983 ( .B1(n386), .B2(n481), .A(n1377), .ZN(n2163) );
  AND2_X4 U984 ( .A1(n331), .A2(n484), .ZN(n1377) );
  XOR2_X2 U985 ( .A(n2130), .B(n289), .Z(n1748) );
  OAI21_X4 U986 ( .B1(n2810), .B2(n3158), .A(n2164), .ZN(n2130) );
  AOI222_X2 U987 ( .A1(n3134), .A2(n484), .B1(n331), .B2(n481), .C1(n386), 
        .C2(n478), .ZN(n2164) );
  XOR2_X2 U988 ( .A(n2131), .B(n289), .Z(n1749) );
  OAI21_X4 U989 ( .B1(n2811), .B2(n3158), .A(n2165), .ZN(n2131) );
  AOI222_X2 U990 ( .A1(n3133), .A2(n481), .B1(n331), .B2(n478), .C1(n386), 
        .C2(n475), .ZN(n2165) );
  XOR2_X2 U991 ( .A(n2132), .B(n289), .Z(n1750) );
  OAI21_X4 U992 ( .B1(n2812), .B2(n3158), .A(n2166), .ZN(n2132) );
  AOI222_X2 U993 ( .A1(n3134), .A2(n478), .B1(n331), .B2(n475), .C1(n386), 
        .C2(n472), .ZN(n2166) );
  XOR2_X2 U994 ( .A(n2133), .B(n289), .Z(n1751) );
  OAI21_X4 U995 ( .B1(n2813), .B2(n3158), .A(n2167), .ZN(n2133) );
  AOI222_X2 U996 ( .A1(n3133), .A2(n475), .B1(n331), .B2(n472), .C1(n386), 
        .C2(n469), .ZN(n2167) );
  XOR2_X2 U997 ( .A(n2134), .B(n289), .Z(n1752) );
  OAI21_X4 U998 ( .B1(n2814), .B2(n3158), .A(n2168), .ZN(n2134) );
  AOI222_X2 U999 ( .A1(n3134), .A2(n472), .B1(n331), .B2(n469), .C1(n386), 
        .C2(n466), .ZN(n2168) );
  XOR2_X2 U1000 ( .A(n2135), .B(n289), .Z(n1753) );
  OAI21_X4 U1001 ( .B1(n2815), .B2(n3158), .A(n2169), .ZN(n2135) );
  AOI222_X2 U1002 ( .A1(n3133), .A2(n469), .B1(n331), .B2(n466), .C1(n386), 
        .C2(n463), .ZN(n2169) );
  XOR2_X2 U1003 ( .A(n2136), .B(n289), .Z(n1754) );
  OAI21_X4 U1004 ( .B1(n2816), .B2(n3158), .A(n2170), .ZN(n2136) );
  AOI222_X2 U1005 ( .A1(n3134), .A2(n466), .B1(n331), .B2(n463), .C1(n386), 
        .C2(n460), .ZN(n2170) );
  XOR2_X2 U1006 ( .A(n2137), .B(n289), .Z(n1755) );
  OAI21_X4 U1007 ( .B1(n2817), .B2(n3158), .A(n2171), .ZN(n2137) );
  AOI222_X2 U1008 ( .A1(n3133), .A2(n463), .B1(n331), .B2(n460), .C1(n386), 
        .C2(n457), .ZN(n2171) );
  XOR2_X2 U1009 ( .A(n2138), .B(n289), .Z(n1756) );
  OAI21_X4 U1010 ( .B1(n2818), .B2(n3158), .A(n2172), .ZN(n2138) );
  AOI222_X2 U1011 ( .A1(n3134), .A2(n460), .B1(n331), .B2(n457), .C1(n386), 
        .C2(n454), .ZN(n2172) );
  XOR2_X2 U1012 ( .A(n2139), .B(n289), .Z(n1757) );
  OAI21_X4 U1013 ( .B1(n2819), .B2(n3158), .A(n2173), .ZN(n2139) );
  AOI222_X2 U1014 ( .A1(n3134), .A2(n457), .B1(n331), .B2(n454), .C1(n386), 
        .C2(n451), .ZN(n2173) );
  XOR2_X2 U1015 ( .A(n2140), .B(n289), .Z(n1758) );
  OAI21_X4 U1016 ( .B1(n2820), .B2(n3158), .A(n2174), .ZN(n2140) );
  AOI222_X2 U1017 ( .A1(n3133), .A2(n454), .B1(n331), .B2(n451), .C1(n386), 
        .C2(n448), .ZN(n2174) );
  XOR2_X2 U1018 ( .A(n2141), .B(n289), .Z(n1759) );
  OAI21_X4 U1019 ( .B1(n2821), .B2(n3158), .A(n2175), .ZN(n2141) );
  AOI222_X2 U1020 ( .A1(n3133), .A2(n451), .B1(n331), .B2(n448), .C1(n386), 
        .C2(n445), .ZN(n2175) );
  XOR2_X2 U1021 ( .A(n2142), .B(n289), .Z(n1760) );
  OAI21_X4 U1022 ( .B1(n2822), .B2(n3158), .A(n2176), .ZN(n2142) );
  AOI222_X2 U1023 ( .A1(n3134), .A2(n448), .B1(n331), .B2(n445), .C1(n386), 
        .C2(n442), .ZN(n2176) );
  XOR2_X2 U1024 ( .A(n2143), .B(n289), .Z(n1761) );
  OAI21_X4 U1025 ( .B1(n2823), .B2(n3158), .A(n2177), .ZN(n2143) );
  AOI222_X2 U1026 ( .A1(n3133), .A2(n445), .B1(n331), .B2(n442), .C1(n386), 
        .C2(n439), .ZN(n2177) );
  XOR2_X2 U1027 ( .A(n2144), .B(n289), .Z(n1762) );
  OAI21_X4 U1028 ( .B1(n2824), .B2(n3158), .A(n2178), .ZN(n2144) );
  AOI222_X2 U1029 ( .A1(n3134), .A2(n442), .B1(n331), .B2(n439), .C1(n386), 
        .C2(n436), .ZN(n2178) );
  XOR2_X2 U1030 ( .A(n2145), .B(n289), .Z(n1763) );
  OAI21_X4 U1031 ( .B1(n2825), .B2(n3158), .A(n2179), .ZN(n2145) );
  AOI222_X2 U1032 ( .A1(n3133), .A2(n439), .B1(n331), .B2(n436), .C1(n386), 
        .C2(n433), .ZN(n2179) );
  XOR2_X2 U1033 ( .A(n2146), .B(n289), .Z(n1764) );
  OAI21_X4 U1034 ( .B1(n2826), .B2(n3158), .A(n2180), .ZN(n2146) );
  AOI222_X2 U1035 ( .A1(n3134), .A2(n436), .B1(n331), .B2(n433), .C1(n386), 
        .C2(n430), .ZN(n2180) );
  XOR2_X2 U1036 ( .A(n2147), .B(n289), .Z(n907) );
  OAI21_X4 U1037 ( .B1(n2827), .B2(n3158), .A(n2181), .ZN(n2147) );
  AOI222_X2 U1038 ( .A1(n3133), .A2(n433), .B1(n331), .B2(n430), .C1(n386), 
        .C2(n427), .ZN(n2181) );
  XOR2_X2 U1039 ( .A(n2148), .B(n289), .Z(n1765) );
  OAI21_X4 U1040 ( .B1(n2828), .B2(n3158), .A(n2182), .ZN(n2148) );
  AOI222_X2 U1041 ( .A1(n3134), .A2(n430), .B1(n331), .B2(n427), .C1(n386), 
        .C2(n424), .ZN(n2182) );
  XOR2_X2 U1042 ( .A(n2149), .B(n289), .Z(n1766) );
  OAI21_X4 U1043 ( .B1(n2829), .B2(n3158), .A(n2183), .ZN(n2149) );
  AOI222_X2 U1044 ( .A1(n3133), .A2(n427), .B1(n331), .B2(n424), .C1(n386), 
        .C2(n421), .ZN(n2183) );
  XOR2_X2 U1045 ( .A(n2150), .B(n289), .Z(n1767) );
  OAI21_X4 U1046 ( .B1(n2830), .B2(n3158), .A(n2184), .ZN(n2150) );
  AOI222_X2 U1047 ( .A1(n3134), .A2(n424), .B1(n331), .B2(n421), .C1(n386), 
        .C2(n418), .ZN(n2184) );
  XOR2_X2 U1048 ( .A(n2151), .B(n289), .Z(n1768) );
  OAI21_X4 U1049 ( .B1(n2831), .B2(n3158), .A(n2185), .ZN(n2151) );
  AOI222_X2 U1050 ( .A1(n3133), .A2(n421), .B1(n331), .B2(n418), .C1(n386), 
        .C2(n415), .ZN(n2185) );
  XOR2_X2 U1051 ( .A(n2152), .B(n289), .Z(n1769) );
  OAI21_X4 U1052 ( .B1(n2832), .B2(n3158), .A(n2186), .ZN(n2152) );
  AOI222_X2 U1053 ( .A1(n3134), .A2(n418), .B1(n331), .B2(n415), .C1(n386), 
        .C2(n412), .ZN(n2186) );
  XOR2_X2 U1054 ( .A(n2153), .B(n289), .Z(n1770) );
  OAI21_X4 U1055 ( .B1(n2833), .B2(n3158), .A(n2187), .ZN(n2153) );
  AOI222_X2 U1056 ( .A1(n3133), .A2(n415), .B1(n331), .B2(n412), .C1(n386), 
        .C2(n409), .ZN(n2187) );
  XOR2_X2 U1057 ( .A(n2154), .B(n289), .Z(n1771) );
  OAI21_X4 U1058 ( .B1(n2834), .B2(n3157), .A(n2188), .ZN(n2154) );
  AOI222_X2 U1059 ( .A1(n3134), .A2(n412), .B1(n331), .B2(n409), .C1(n386), 
        .C2(n406), .ZN(n2188) );
  XOR2_X2 U1060 ( .A(n2155), .B(n289), .Z(n1772) );
  OAI21_X4 U1061 ( .B1(n2835), .B2(n3157), .A(n2189), .ZN(n2155) );
  AOI222_X2 U1062 ( .A1(n3133), .A2(n409), .B1(n331), .B2(n406), .C1(n386), 
        .C2(n403), .ZN(n2189) );
  XOR2_X2 U1063 ( .A(n2156), .B(n289), .Z(n1773) );
  OAI21_X4 U1064 ( .B1(n2836), .B2(n3157), .A(n2190), .ZN(n2156) );
  AOI222_X2 U1065 ( .A1(n3134), .A2(n406), .B1(n331), .B2(n403), .C1(n386), 
        .C2(n400), .ZN(n2190) );
  XOR2_X2 U1066 ( .A(n2157), .B(n289), .Z(n1774) );
  OAI21_X4 U1067 ( .B1(n2837), .B2(n3157), .A(n2191), .ZN(n2157) );
  AOI222_X2 U1068 ( .A1(n3133), .A2(n403), .B1(n331), .B2(n400), .C1(n386), 
        .C2(n397), .ZN(n2191) );
  XOR2_X2 U1069 ( .A(n2158), .B(n289), .Z(n1775) );
  OAI21_X4 U1070 ( .B1(n2838), .B2(n3157), .A(n2192), .ZN(n2158) );
  AOI222_X2 U1071 ( .A1(n3134), .A2(n400), .B1(n331), .B2(n397), .C1(n386), 
        .C2(n393), .ZN(n2192) );
  XOR2_X2 U1072 ( .A(n2159), .B(n289), .Z(n1776) );
  OAI21_X4 U1073 ( .B1(n2839), .B2(n3157), .A(n2193), .ZN(n2159) );
  AOI222_X2 U1074 ( .A1(n3133), .A2(n397), .B1(n331), .B2(n393), .C1(n386), 
        .C2(n390), .ZN(n2193) );
  XOR2_X2 U1075 ( .A(n2160), .B(n289), .Z(n1777) );
  OAI21_X4 U1076 ( .B1(n2840), .B2(n3157), .A(n2194), .ZN(n2160) );
  XOR2_X2 U1078 ( .A(n2161), .B(n289), .Z(n1778) );
  OAI21_X4 U1079 ( .B1(n2841), .B2(n3157), .A(n2195), .ZN(n2161) );
  AND2_X4 U1081 ( .A1(n3133), .A2(n390), .ZN(n1379) );
  XOR2_X2 U1083 ( .A(n2196), .B(n286), .Z(n1780) );
  OAI21_X4 U1084 ( .B1(n2808), .B2(n3155), .A(n2230), .ZN(n2196) );
  NAND2_X4 U1085 ( .A1(n384), .A2(n484), .ZN(n2230) );
  XOR2_X2 U1086 ( .A(n2197), .B(n286), .Z(n1781) );
  OAI21_X4 U1087 ( .B1(n2809), .B2(n3155), .A(n2231), .ZN(n2197) );
  AOI21_X4 U1088 ( .B1(n384), .B2(n481), .A(n1380), .ZN(n2231) );
  AND2_X4 U1089 ( .A1(n329), .A2(n484), .ZN(n1380) );
  XOR2_X2 U1090 ( .A(n2198), .B(n286), .Z(n1782) );
  OAI21_X4 U1091 ( .B1(n2810), .B2(n3155), .A(n2232), .ZN(n2198) );
  AOI222_X2 U1092 ( .A1(n3137), .A2(n484), .B1(n329), .B2(n481), .C1(n384), 
        .C2(n478), .ZN(n2232) );
  XOR2_X2 U1093 ( .A(n2199), .B(n286), .Z(n1783) );
  OAI21_X4 U1094 ( .B1(n2811), .B2(n3155), .A(n2233), .ZN(n2199) );
  AOI222_X2 U1095 ( .A1(n3136), .A2(n481), .B1(n329), .B2(n478), .C1(n384), 
        .C2(n475), .ZN(n2233) );
  XOR2_X2 U1096 ( .A(n2200), .B(n286), .Z(n1784) );
  OAI21_X4 U1097 ( .B1(n2812), .B2(n3155), .A(n2234), .ZN(n2200) );
  AOI222_X2 U1098 ( .A1(n3137), .A2(n478), .B1(n329), .B2(n475), .C1(n384), 
        .C2(n472), .ZN(n2234) );
  XOR2_X2 U1099 ( .A(n2201), .B(n286), .Z(n1785) );
  OAI21_X4 U1100 ( .B1(n2813), .B2(n3155), .A(n2235), .ZN(n2201) );
  AOI222_X2 U1101 ( .A1(n3136), .A2(n475), .B1(n329), .B2(n472), .C1(n384), 
        .C2(n469), .ZN(n2235) );
  XOR2_X2 U1102 ( .A(n2202), .B(n286), .Z(n1786) );
  OAI21_X4 U1103 ( .B1(n2814), .B2(n3155), .A(n2236), .ZN(n2202) );
  AOI222_X2 U1104 ( .A1(n3137), .A2(n472), .B1(n329), .B2(n469), .C1(n384), 
        .C2(n466), .ZN(n2236) );
  XOR2_X2 U1105 ( .A(n2203), .B(n286), .Z(n1787) );
  OAI21_X4 U1106 ( .B1(n2815), .B2(n3155), .A(n2237), .ZN(n2203) );
  AOI222_X2 U1107 ( .A1(n3136), .A2(n469), .B1(n329), .B2(n466), .C1(n384), 
        .C2(n463), .ZN(n2237) );
  XOR2_X2 U1108 ( .A(n2204), .B(n286), .Z(n1788) );
  OAI21_X4 U1109 ( .B1(n2816), .B2(n3155), .A(n2238), .ZN(n2204) );
  AOI222_X2 U1110 ( .A1(n3137), .A2(n466), .B1(n329), .B2(n463), .C1(n384), 
        .C2(n460), .ZN(n2238) );
  XOR2_X2 U1111 ( .A(n2205), .B(n286), .Z(n1789) );
  OAI21_X4 U1112 ( .B1(n2817), .B2(n3155), .A(n2239), .ZN(n2205) );
  AOI222_X2 U1113 ( .A1(n3136), .A2(n463), .B1(n329), .B2(n460), .C1(n384), 
        .C2(n457), .ZN(n2239) );
  XOR2_X2 U1114 ( .A(n2206), .B(n286), .Z(n1790) );
  OAI21_X4 U1115 ( .B1(n2818), .B2(n3155), .A(n2240), .ZN(n2206) );
  AOI222_X2 U1116 ( .A1(n3137), .A2(n460), .B1(n329), .B2(n457), .C1(n384), 
        .C2(n454), .ZN(n2240) );
  XOR2_X2 U1117 ( .A(n2207), .B(n286), .Z(n1791) );
  OAI21_X4 U1118 ( .B1(n2819), .B2(n3155), .A(n2241), .ZN(n2207) );
  AOI222_X2 U1119 ( .A1(n3136), .A2(n457), .B1(n329), .B2(n454), .C1(n384), 
        .C2(n451), .ZN(n2241) );
  XOR2_X2 U1120 ( .A(n2208), .B(n286), .Z(n1792) );
  OAI21_X4 U1121 ( .B1(n2820), .B2(n3155), .A(n2242), .ZN(n2208) );
  AOI222_X2 U1122 ( .A1(n3137), .A2(n454), .B1(n329), .B2(n451), .C1(n384), 
        .C2(n448), .ZN(n2242) );
  XOR2_X2 U1123 ( .A(n2209), .B(n286), .Z(n1793) );
  OAI21_X4 U1124 ( .B1(n2821), .B2(n3155), .A(n2243), .ZN(n2209) );
  AOI222_X2 U1125 ( .A1(n3136), .A2(n451), .B1(n329), .B2(n448), .C1(n384), 
        .C2(n445), .ZN(n2243) );
  XOR2_X2 U1126 ( .A(n2210), .B(n286), .Z(n1794) );
  OAI21_X4 U1127 ( .B1(n2822), .B2(n3155), .A(n2244), .ZN(n2210) );
  AOI222_X2 U1128 ( .A1(n3137), .A2(n448), .B1(n329), .B2(n445), .C1(n384), 
        .C2(n442), .ZN(n2244) );
  XOR2_X2 U1129 ( .A(n2211), .B(n286), .Z(n1795) );
  OAI21_X4 U1130 ( .B1(n2823), .B2(n3155), .A(n2245), .ZN(n2211) );
  AOI222_X2 U1131 ( .A1(n3136), .A2(n445), .B1(n329), .B2(n442), .C1(n384), 
        .C2(n439), .ZN(n2245) );
  XOR2_X2 U1132 ( .A(n2212), .B(n286), .Z(n1796) );
  OAI21_X4 U1133 ( .B1(n2824), .B2(n3155), .A(n2246), .ZN(n2212) );
  AOI222_X2 U1134 ( .A1(n3137), .A2(n442), .B1(n329), .B2(n439), .C1(n384), 
        .C2(n436), .ZN(n2246) );
  XOR2_X2 U1135 ( .A(n2213), .B(n286), .Z(n1797) );
  OAI21_X4 U1136 ( .B1(n2825), .B2(n3155), .A(n2247), .ZN(n2213) );
  AOI222_X2 U1137 ( .A1(n3136), .A2(n439), .B1(n329), .B2(n436), .C1(n384), 
        .C2(n433), .ZN(n2247) );
  XOR2_X2 U1138 ( .A(n2214), .B(n286), .Z(n1798) );
  OAI21_X4 U1139 ( .B1(n2826), .B2(n3155), .A(n2248), .ZN(n2214) );
  AOI222_X2 U1140 ( .A1(n3137), .A2(n436), .B1(n329), .B2(n433), .C1(n384), 
        .C2(n430), .ZN(n2248) );
  XOR2_X2 U1141 ( .A(n2215), .B(n286), .Z(n1799) );
  OAI21_X4 U1142 ( .B1(n2827), .B2(n3155), .A(n2249), .ZN(n2215) );
  AOI222_X2 U1143 ( .A1(n3136), .A2(n433), .B1(n329), .B2(n430), .C1(n384), 
        .C2(n427), .ZN(n2249) );
  XOR2_X2 U1144 ( .A(n2216), .B(n286), .Z(n1800) );
  OAI21_X4 U1145 ( .B1(n2828), .B2(n3155), .A(n2250), .ZN(n2216) );
  AOI222_X2 U1146 ( .A1(n3137), .A2(n430), .B1(n329), .B2(n427), .C1(n384), 
        .C2(n424), .ZN(n2250) );
  XOR2_X2 U1147 ( .A(n2217), .B(n286), .Z(n1801) );
  OAI21_X4 U1148 ( .B1(n2829), .B2(n3155), .A(n2251), .ZN(n2217) );
  AOI222_X2 U1149 ( .A1(n3136), .A2(n427), .B1(n329), .B2(n424), .C1(n384), 
        .C2(n421), .ZN(n2251) );
  XOR2_X2 U1150 ( .A(n2218), .B(n286), .Z(n1802) );
  OAI21_X4 U1151 ( .B1(n2830), .B2(n3155), .A(n2252), .ZN(n2218) );
  AOI222_X2 U1152 ( .A1(n3137), .A2(n424), .B1(n329), .B2(n421), .C1(n384), 
        .C2(n418), .ZN(n2252) );
  XOR2_X2 U1153 ( .A(n2219), .B(n286), .Z(n1803) );
  OAI21_X4 U1154 ( .B1(n2831), .B2(n3155), .A(n2253), .ZN(n2219) );
  AOI222_X2 U1155 ( .A1(n3136), .A2(n421), .B1(n329), .B2(n418), .C1(n384), 
        .C2(n415), .ZN(n2253) );
  XOR2_X2 U1156 ( .A(n2220), .B(n286), .Z(n1804) );
  OAI21_X4 U1157 ( .B1(n2832), .B2(n3155), .A(n2254), .ZN(n2220) );
  AOI222_X2 U1158 ( .A1(n3137), .A2(n418), .B1(n329), .B2(n415), .C1(n384), 
        .C2(n412), .ZN(n2254) );
  XOR2_X2 U1159 ( .A(n2221), .B(n286), .Z(n1805) );
  OAI21_X4 U1160 ( .B1(n2833), .B2(n3155), .A(n2255), .ZN(n2221) );
  AOI222_X2 U1161 ( .A1(n3136), .A2(n415), .B1(n329), .B2(n412), .C1(n384), 
        .C2(n409), .ZN(n2255) );
  XOR2_X2 U1162 ( .A(n2222), .B(n286), .Z(n1806) );
  OAI21_X4 U1163 ( .B1(n2834), .B2(n3154), .A(n2256), .ZN(n2222) );
  AOI222_X2 U1164 ( .A1(n3137), .A2(n412), .B1(n329), .B2(n409), .C1(n384), 
        .C2(n406), .ZN(n2256) );
  XOR2_X2 U1165 ( .A(n2223), .B(n286), .Z(n1807) );
  OAI21_X4 U1166 ( .B1(n2835), .B2(n3154), .A(n2257), .ZN(n2223) );
  AOI222_X2 U1167 ( .A1(n3136), .A2(n409), .B1(n329), .B2(n406), .C1(n384), 
        .C2(n403), .ZN(n2257) );
  XOR2_X2 U1168 ( .A(n2224), .B(n286), .Z(n1808) );
  OAI21_X4 U1169 ( .B1(n2836), .B2(n3154), .A(n2258), .ZN(n2224) );
  AOI222_X2 U1170 ( .A1(n3137), .A2(n406), .B1(n329), .B2(n403), .C1(n384), 
        .C2(n400), .ZN(n2258) );
  XOR2_X2 U1171 ( .A(n2225), .B(n286), .Z(n1809) );
  OAI21_X4 U1172 ( .B1(n2837), .B2(n3154), .A(n2259), .ZN(n2225) );
  AOI222_X2 U1173 ( .A1(n3136), .A2(n403), .B1(n329), .B2(n400), .C1(n384), 
        .C2(n397), .ZN(n2259) );
  XOR2_X2 U1174 ( .A(n2226), .B(n286), .Z(n1810) );
  OAI21_X4 U1175 ( .B1(n2838), .B2(n3154), .A(n2260), .ZN(n2226) );
  AOI222_X2 U1176 ( .A1(n3137), .A2(n400), .B1(n329), .B2(n397), .C1(n384), 
        .C2(n393), .ZN(n2260) );
  XOR2_X2 U1177 ( .A(n2227), .B(n286), .Z(n1811) );
  OAI21_X4 U1178 ( .B1(n2839), .B2(n3154), .A(n2261), .ZN(n2227) );
  AOI222_X2 U1179 ( .A1(n3136), .A2(n397), .B1(n329), .B2(n393), .C1(n384), 
        .C2(n390), .ZN(n2261) );
  XOR2_X2 U1180 ( .A(n2228), .B(n286), .Z(n1812) );
  OAI21_X4 U1181 ( .B1(n2840), .B2(n3154), .A(n2262), .ZN(n2228) );
  XOR2_X2 U1183 ( .A(n2229), .B(n286), .Z(n1813) );
  OAI21_X4 U1184 ( .B1(n2841), .B2(n3154), .A(n2263), .ZN(n2229) );
  AND2_X4 U1186 ( .A1(n3136), .A2(n390), .ZN(n1382) );
  XOR2_X2 U1188 ( .A(n2264), .B(n283), .Z(n1815) );
  OAI21_X4 U1189 ( .B1(n2808), .B2(n3162), .A(n2298), .ZN(n2264) );
  NAND2_X4 U1190 ( .A1(n382), .A2(n484), .ZN(n2298) );
  XOR2_X2 U1191 ( .A(n2265), .B(n283), .Z(n1816) );
  OAI21_X4 U1192 ( .B1(n2809), .B2(n3162), .A(n2299), .ZN(n2265) );
  AOI21_X4 U1193 ( .B1(n382), .B2(n481), .A(n1383), .ZN(n2299) );
  AND2_X4 U1194 ( .A1(n327), .A2(n484), .ZN(n1383) );
  XOR2_X2 U1195 ( .A(n2266), .B(n283), .Z(n1817) );
  OAI21_X4 U1196 ( .B1(n2810), .B2(n357), .A(n2300), .ZN(n2266) );
  AOI222_X2 U1197 ( .A1(n3140), .A2(n484), .B1(n327), .B2(n481), .C1(n382), 
        .C2(n478), .ZN(n2300) );
  XOR2_X2 U1198 ( .A(n2267), .B(n283), .Z(n1818) );
  OAI21_X4 U1199 ( .B1(n2811), .B2(n357), .A(n2301), .ZN(n2267) );
  AOI222_X2 U1200 ( .A1(n3139), .A2(n481), .B1(n327), .B2(n478), .C1(n382), 
        .C2(n475), .ZN(n2301) );
  XOR2_X2 U1201 ( .A(n2268), .B(n283), .Z(n1819) );
  OAI21_X4 U1202 ( .B1(n2812), .B2(n357), .A(n2302), .ZN(n2268) );
  AOI222_X2 U1203 ( .A1(n3140), .A2(n478), .B1(n327), .B2(n475), .C1(n382), 
        .C2(n472), .ZN(n2302) );
  XOR2_X2 U1204 ( .A(n2269), .B(n283), .Z(n1820) );
  OAI21_X4 U1205 ( .B1(n2813), .B2(n357), .A(n2303), .ZN(n2269) );
  AOI222_X2 U1206 ( .A1(n3139), .A2(n475), .B1(n327), .B2(n472), .C1(n382), 
        .C2(n469), .ZN(n2303) );
  XOR2_X2 U1207 ( .A(n2270), .B(n283), .Z(n1821) );
  OAI21_X4 U1208 ( .B1(n2814), .B2(n357), .A(n2304), .ZN(n2270) );
  AOI222_X2 U1209 ( .A1(n3140), .A2(n472), .B1(n327), .B2(n469), .C1(n382), 
        .C2(n466), .ZN(n2304) );
  XOR2_X2 U1210 ( .A(n2271), .B(n283), .Z(n1822) );
  OAI21_X4 U1211 ( .B1(n2815), .B2(n357), .A(n2305), .ZN(n2271) );
  AOI222_X2 U1212 ( .A1(n3139), .A2(n469), .B1(n327), .B2(n466), .C1(n382), 
        .C2(n463), .ZN(n2305) );
  XOR2_X2 U1213 ( .A(n2272), .B(n283), .Z(n1823) );
  OAI21_X4 U1214 ( .B1(n2816), .B2(n357), .A(n2306), .ZN(n2272) );
  AOI222_X2 U1215 ( .A1(n3140), .A2(n466), .B1(n327), .B2(n463), .C1(n382), 
        .C2(n460), .ZN(n2306) );
  XOR2_X2 U1216 ( .A(n2273), .B(n283), .Z(n1824) );
  OAI21_X4 U1217 ( .B1(n2817), .B2(n357), .A(n2307), .ZN(n2273) );
  AOI222_X2 U1218 ( .A1(n3139), .A2(n463), .B1(n327), .B2(n460), .C1(n382), 
        .C2(n457), .ZN(n2307) );
  XOR2_X2 U1219 ( .A(n2274), .B(n283), .Z(n1825) );
  OAI21_X4 U1220 ( .B1(n2818), .B2(n357), .A(n2308), .ZN(n2274) );
  AOI222_X2 U1221 ( .A1(n3140), .A2(n460), .B1(n327), .B2(n457), .C1(n382), 
        .C2(n454), .ZN(n2308) );
  XOR2_X2 U1222 ( .A(n2275), .B(n283), .Z(n1826) );
  OAI21_X4 U1223 ( .B1(n2819), .B2(n357), .A(n2309), .ZN(n2275) );
  AOI222_X2 U1224 ( .A1(n3139), .A2(n457), .B1(n327), .B2(n454), .C1(n382), 
        .C2(n451), .ZN(n2309) );
  XOR2_X2 U1225 ( .A(n2276), .B(n283), .Z(n1827) );
  OAI21_X4 U1226 ( .B1(n2820), .B2(n357), .A(n2310), .ZN(n2276) );
  AOI222_X2 U1227 ( .A1(n3140), .A2(n454), .B1(n327), .B2(n451), .C1(n382), 
        .C2(n448), .ZN(n2310) );
  XOR2_X2 U1228 ( .A(n2277), .B(n283), .Z(n1828) );
  OAI21_X4 U1229 ( .B1(n2821), .B2(n357), .A(n2311), .ZN(n2277) );
  AOI222_X2 U1230 ( .A1(n3139), .A2(n451), .B1(n327), .B2(n448), .C1(n382), 
        .C2(n445), .ZN(n2311) );
  XOR2_X2 U1231 ( .A(n2278), .B(n283), .Z(n1829) );
  OAI21_X4 U1232 ( .B1(n2822), .B2(n357), .A(n2312), .ZN(n2278) );
  AOI222_X2 U1233 ( .A1(n3140), .A2(n448), .B1(n327), .B2(n445), .C1(n382), 
        .C2(n442), .ZN(n2312) );
  XOR2_X2 U1234 ( .A(n2279), .B(n283), .Z(n1830) );
  OAI21_X4 U1235 ( .B1(n2823), .B2(n357), .A(n2313), .ZN(n2279) );
  AOI222_X2 U1236 ( .A1(n3139), .A2(n445), .B1(n327), .B2(n442), .C1(n382), 
        .C2(n439), .ZN(n2313) );
  XOR2_X2 U1237 ( .A(n2280), .B(n283), .Z(n1831) );
  OAI21_X4 U1238 ( .B1(n2824), .B2(n357), .A(n2314), .ZN(n2280) );
  AOI222_X2 U1239 ( .A1(n3140), .A2(n442), .B1(n327), .B2(n439), .C1(n382), 
        .C2(n436), .ZN(n2314) );
  XOR2_X2 U1240 ( .A(n2281), .B(n283), .Z(n1832) );
  OAI21_X4 U1241 ( .B1(n2825), .B2(n357), .A(n2315), .ZN(n2281) );
  AOI222_X2 U1242 ( .A1(n3139), .A2(n439), .B1(n327), .B2(n436), .C1(n382), 
        .C2(n433), .ZN(n2315) );
  XOR2_X2 U1243 ( .A(n2282), .B(n283), .Z(n1833) );
  OAI21_X4 U1244 ( .B1(n2826), .B2(n357), .A(n2316), .ZN(n2282) );
  AOI222_X2 U1245 ( .A1(n3140), .A2(n436), .B1(n327), .B2(n433), .C1(n382), 
        .C2(n430), .ZN(n2316) );
  XOR2_X2 U1246 ( .A(n2283), .B(n283), .Z(n1834) );
  OAI21_X4 U1247 ( .B1(n2827), .B2(n357), .A(n2317), .ZN(n2283) );
  AOI222_X2 U1248 ( .A1(n3139), .A2(n433), .B1(n327), .B2(n430), .C1(n382), 
        .C2(n427), .ZN(n2317) );
  XOR2_X2 U1249 ( .A(n2284), .B(n283), .Z(n1835) );
  OAI21_X4 U1250 ( .B1(n2828), .B2(n357), .A(n2318), .ZN(n2284) );
  AOI222_X2 U1251 ( .A1(n3140), .A2(n430), .B1(n327), .B2(n427), .C1(n382), 
        .C2(n424), .ZN(n2318) );
  XOR2_X2 U1252 ( .A(n2285), .B(n283), .Z(n1836) );
  OAI21_X4 U1253 ( .B1(n2829), .B2(n357), .A(n2319), .ZN(n2285) );
  AOI222_X2 U1254 ( .A1(n3140), .A2(n427), .B1(n327), .B2(n424), .C1(n382), 
        .C2(n421), .ZN(n2319) );
  XOR2_X2 U1255 ( .A(n2286), .B(n283), .Z(n1837) );
  OAI21_X4 U1256 ( .B1(n2830), .B2(n357), .A(n2320), .ZN(n2286) );
  AOI222_X2 U1257 ( .A1(n3139), .A2(n424), .B1(n327), .B2(n421), .C1(n382), 
        .C2(n418), .ZN(n2320) );
  XOR2_X2 U1258 ( .A(n2287), .B(n283), .Z(n1838) );
  OAI21_X4 U1259 ( .B1(n2831), .B2(n357), .A(n2321), .ZN(n2287) );
  AOI222_X2 U1260 ( .A1(n3139), .A2(n421), .B1(n327), .B2(n418), .C1(n382), 
        .C2(n415), .ZN(n2321) );
  XOR2_X2 U1261 ( .A(n2288), .B(n283), .Z(n1839) );
  OAI21_X4 U1262 ( .B1(n2832), .B2(n357), .A(n2322), .ZN(n2288) );
  AOI222_X2 U1263 ( .A1(n3139), .A2(n418), .B1(n327), .B2(n415), .C1(n382), 
        .C2(n412), .ZN(n2322) );
  XOR2_X2 U1264 ( .A(n2289), .B(n283), .Z(n1840) );
  OAI21_X4 U1265 ( .B1(n2833), .B2(n357), .A(n2323), .ZN(n2289) );
  AOI222_X2 U1266 ( .A1(n3140), .A2(n415), .B1(n327), .B2(n412), .C1(n382), 
        .C2(n409), .ZN(n2323) );
  XOR2_X2 U1267 ( .A(n2290), .B(n283), .Z(n1841) );
  OAI21_X4 U1268 ( .B1(n2834), .B2(n357), .A(n2324), .ZN(n2290) );
  AOI222_X2 U1269 ( .A1(n3140), .A2(n412), .B1(n327), .B2(n409), .C1(n382), 
        .C2(n406), .ZN(n2324) );
  XOR2_X2 U1270 ( .A(n2291), .B(n283), .Z(n1842) );
  OAI21_X4 U1271 ( .B1(n2835), .B2(n357), .A(n2325), .ZN(n2291) );
  AOI222_X2 U1272 ( .A1(n3140), .A2(n409), .B1(n327), .B2(n406), .C1(n382), 
        .C2(n403), .ZN(n2325) );
  XOR2_X2 U1273 ( .A(n2292), .B(n283), .Z(n1843) );
  OAI21_X4 U1274 ( .B1(n2836), .B2(n357), .A(n2326), .ZN(n2292) );
  AOI222_X2 U1275 ( .A1(n3139), .A2(n406), .B1(n327), .B2(n403), .C1(n382), 
        .C2(n400), .ZN(n2326) );
  XOR2_X2 U1276 ( .A(n2293), .B(n283), .Z(n1844) );
  OAI21_X4 U1277 ( .B1(n2837), .B2(n357), .A(n2327), .ZN(n2293) );
  AOI222_X2 U1278 ( .A1(n3139), .A2(n403), .B1(n327), .B2(n400), .C1(n382), 
        .C2(n397), .ZN(n2327) );
  XOR2_X2 U1279 ( .A(n2294), .B(n283), .Z(n1845) );
  OAI21_X4 U1280 ( .B1(n2838), .B2(n357), .A(n2328), .ZN(n2294) );
  AOI222_X2 U1281 ( .A1(n3140), .A2(n400), .B1(n327), .B2(n397), .C1(n382), 
        .C2(n393), .ZN(n2328) );
  XOR2_X2 U1282 ( .A(n2295), .B(n283), .Z(n1846) );
  OAI21_X4 U1283 ( .B1(n2839), .B2(n357), .A(n2329), .ZN(n2295) );
  AOI222_X2 U1284 ( .A1(n3139), .A2(n397), .B1(n327), .B2(n393), .C1(n382), 
        .C2(n390), .ZN(n2329) );
  XOR2_X2 U1285 ( .A(n2296), .B(n283), .Z(n1847) );
  OAI21_X4 U1286 ( .B1(n2840), .B2(n357), .A(n2330), .ZN(n2296) );
  XOR2_X2 U1288 ( .A(n2297), .B(n283), .Z(n1848) );
  OAI21_X4 U1289 ( .B1(n2841), .B2(n357), .A(n2331), .ZN(n2297) );
  AND2_X4 U1291 ( .A1(n3139), .A2(n390), .ZN(n1385) );
  XOR2_X2 U1293 ( .A(n2332), .B(n280), .Z(n1850) );
  OAI21_X4 U1294 ( .B1(n2808), .B2(n3128), .A(n2366), .ZN(n2332) );
  NAND2_X4 U1295 ( .A1(n380), .A2(n484), .ZN(n2366) );
  XOR2_X2 U1296 ( .A(n2333), .B(n280), .Z(n1851) );
  OAI21_X4 U1297 ( .B1(n2809), .B2(n3128), .A(n2367), .ZN(n2333) );
  AOI21_X4 U1298 ( .B1(n380), .B2(n481), .A(n1386), .ZN(n2367) );
  AND2_X4 U1299 ( .A1(n325), .A2(n484), .ZN(n1386) );
  XOR2_X2 U1300 ( .A(n2334), .B(n280), .Z(n1852) );
  OAI21_X4 U1301 ( .B1(n2810), .B2(n354), .A(n2368), .ZN(n2334) );
  AOI222_X2 U1302 ( .A1(n3143), .A2(n484), .B1(n325), .B2(n481), .C1(n380), 
        .C2(n478), .ZN(n2368) );
  XOR2_X2 U1303 ( .A(n2335), .B(n280), .Z(n1853) );
  OAI21_X4 U1304 ( .B1(n2811), .B2(n354), .A(n2369), .ZN(n2335) );
  AOI222_X2 U1305 ( .A1(n3142), .A2(n481), .B1(n325), .B2(n478), .C1(n380), 
        .C2(n475), .ZN(n2369) );
  XOR2_X2 U1306 ( .A(n2336), .B(n280), .Z(n1854) );
  OAI21_X4 U1307 ( .B1(n2812), .B2(n354), .A(n2370), .ZN(n2336) );
  AOI222_X2 U1308 ( .A1(n3143), .A2(n478), .B1(n325), .B2(n475), .C1(n380), 
        .C2(n472), .ZN(n2370) );
  XOR2_X2 U1309 ( .A(n2337), .B(n280), .Z(n1855) );
  OAI21_X4 U1310 ( .B1(n2813), .B2(n354), .A(n2371), .ZN(n2337) );
  AOI222_X2 U1311 ( .A1(n3142), .A2(n475), .B1(n325), .B2(n472), .C1(n380), 
        .C2(n469), .ZN(n2371) );
  XOR2_X2 U1312 ( .A(n2338), .B(n280), .Z(n1856) );
  OAI21_X4 U1313 ( .B1(n2814), .B2(n354), .A(n2372), .ZN(n2338) );
  AOI222_X2 U1314 ( .A1(n3143), .A2(n472), .B1(n325), .B2(n469), .C1(n380), 
        .C2(n466), .ZN(n2372) );
  XOR2_X2 U1315 ( .A(n2339), .B(n280), .Z(n1857) );
  OAI21_X4 U1316 ( .B1(n2815), .B2(n354), .A(n2373), .ZN(n2339) );
  AOI222_X2 U1317 ( .A1(n3142), .A2(n469), .B1(n325), .B2(n466), .C1(n380), 
        .C2(n463), .ZN(n2373) );
  XOR2_X2 U1318 ( .A(n2340), .B(n280), .Z(n1858) );
  OAI21_X4 U1319 ( .B1(n2816), .B2(n354), .A(n2374), .ZN(n2340) );
  AOI222_X2 U1320 ( .A1(n3143), .A2(n466), .B1(n325), .B2(n463), .C1(n380), 
        .C2(n460), .ZN(n2374) );
  XOR2_X2 U1321 ( .A(n2341), .B(n280), .Z(n1859) );
  OAI21_X4 U1322 ( .B1(n2817), .B2(n354), .A(n2375), .ZN(n2341) );
  AOI222_X2 U1323 ( .A1(n3142), .A2(n463), .B1(n325), .B2(n460), .C1(n380), 
        .C2(n457), .ZN(n2375) );
  XOR2_X2 U1324 ( .A(n2342), .B(n280), .Z(n1860) );
  OAI21_X4 U1325 ( .B1(n2818), .B2(n354), .A(n2376), .ZN(n2342) );
  AOI222_X2 U1326 ( .A1(n3143), .A2(n460), .B1(n325), .B2(n457), .C1(n380), 
        .C2(n454), .ZN(n2376) );
  XOR2_X2 U1327 ( .A(n2343), .B(n280), .Z(n1861) );
  OAI21_X4 U1328 ( .B1(n2819), .B2(n354), .A(n2377), .ZN(n2343) );
  AOI222_X2 U1329 ( .A1(n3142), .A2(n457), .B1(n325), .B2(n454), .C1(n380), 
        .C2(n451), .ZN(n2377) );
  XOR2_X2 U1330 ( .A(n2344), .B(n280), .Z(n1862) );
  OAI21_X4 U1331 ( .B1(n2820), .B2(n354), .A(n2378), .ZN(n2344) );
  AOI222_X2 U1332 ( .A1(n3143), .A2(n454), .B1(n325), .B2(n451), .C1(n380), 
        .C2(n448), .ZN(n2378) );
  XOR2_X2 U1333 ( .A(n2345), .B(n280), .Z(n1863) );
  OAI21_X4 U1334 ( .B1(n2821), .B2(n354), .A(n2379), .ZN(n2345) );
  AOI222_X2 U1335 ( .A1(n3142), .A2(n451), .B1(n325), .B2(n448), .C1(n380), 
        .C2(n445), .ZN(n2379) );
  XOR2_X2 U1336 ( .A(n2346), .B(n280), .Z(n1864) );
  OAI21_X4 U1337 ( .B1(n2822), .B2(n354), .A(n2380), .ZN(n2346) );
  AOI222_X2 U1338 ( .A1(n3142), .A2(n448), .B1(n325), .B2(n445), .C1(n380), 
        .C2(n442), .ZN(n2380) );
  XOR2_X2 U1339 ( .A(n2347), .B(n280), .Z(n1865) );
  OAI21_X4 U1340 ( .B1(n2823), .B2(n354), .A(n2381), .ZN(n2347) );
  AOI222_X2 U1341 ( .A1(n3143), .A2(n445), .B1(n325), .B2(n442), .C1(n380), 
        .C2(n439), .ZN(n2381) );
  XOR2_X2 U1342 ( .A(n2348), .B(n280), .Z(n1866) );
  OAI21_X4 U1343 ( .B1(n2824), .B2(n354), .A(n2382), .ZN(n2348) );
  AOI222_X2 U1344 ( .A1(n3143), .A2(n442), .B1(n325), .B2(n439), .C1(n380), 
        .C2(n436), .ZN(n2382) );
  XOR2_X2 U1345 ( .A(n2349), .B(n280), .Z(n1867) );
  OAI21_X4 U1346 ( .B1(n2825), .B2(n354), .A(n2383), .ZN(n2349) );
  AOI222_X2 U1347 ( .A1(n3142), .A2(n439), .B1(n325), .B2(n436), .C1(n380), 
        .C2(n433), .ZN(n2383) );
  XOR2_X2 U1348 ( .A(n2350), .B(n280), .Z(n1868) );
  OAI21_X4 U1349 ( .B1(n2826), .B2(n354), .A(n2384), .ZN(n2350) );
  AOI222_X2 U1350 ( .A1(n3143), .A2(n436), .B1(n325), .B2(n433), .C1(n380), 
        .C2(n430), .ZN(n2384) );
  XOR2_X2 U1351 ( .A(n2351), .B(n280), .Z(n1869) );
  OAI21_X4 U1352 ( .B1(n2827), .B2(n354), .A(n2385), .ZN(n2351) );
  AOI222_X2 U1353 ( .A1(n3142), .A2(n433), .B1(n325), .B2(n430), .C1(n380), 
        .C2(n427), .ZN(n2385) );
  XOR2_X2 U1354 ( .A(n2352), .B(n280), .Z(n1870) );
  OAI21_X4 U1355 ( .B1(n2828), .B2(n354), .A(n2386), .ZN(n2352) );
  AOI222_X2 U1356 ( .A1(n3143), .A2(n430), .B1(n325), .B2(n427), .C1(n380), 
        .C2(n424), .ZN(n2386) );
  XOR2_X2 U1357 ( .A(n2353), .B(n280), .Z(n1871) );
  OAI21_X4 U1358 ( .B1(n2829), .B2(n354), .A(n2387), .ZN(n2353) );
  AOI222_X2 U1359 ( .A1(n3143), .A2(n427), .B1(n325), .B2(n424), .C1(n380), 
        .C2(n421), .ZN(n2387) );
  XOR2_X2 U1360 ( .A(n2354), .B(n280), .Z(n1872) );
  OAI21_X4 U1361 ( .B1(n2830), .B2(n354), .A(n2388), .ZN(n2354) );
  AOI222_X2 U1362 ( .A1(n3142), .A2(n424), .B1(n325), .B2(n421), .C1(n380), 
        .C2(n418), .ZN(n2388) );
  XOR2_X2 U1363 ( .A(n2355), .B(n280), .Z(n1873) );
  OAI21_X4 U1364 ( .B1(n2831), .B2(n354), .A(n2389), .ZN(n2355) );
  AOI222_X2 U1365 ( .A1(n3142), .A2(n421), .B1(n325), .B2(n418), .C1(n380), 
        .C2(n415), .ZN(n2389) );
  XOR2_X2 U1366 ( .A(n2356), .B(n280), .Z(n1874) );
  OAI21_X4 U1367 ( .B1(n2832), .B2(n354), .A(n2390), .ZN(n2356) );
  AOI222_X2 U1368 ( .A1(n3142), .A2(n418), .B1(n325), .B2(n415), .C1(n380), 
        .C2(n412), .ZN(n2390) );
  XOR2_X2 U1369 ( .A(n2357), .B(n280), .Z(n1875) );
  OAI21_X4 U1370 ( .B1(n2833), .B2(n354), .A(n2391), .ZN(n2357) );
  AOI222_X2 U1371 ( .A1(n3143), .A2(n415), .B1(n325), .B2(n412), .C1(n380), 
        .C2(n409), .ZN(n2391) );
  XOR2_X2 U1372 ( .A(n2358), .B(n280), .Z(n1876) );
  OAI21_X4 U1373 ( .B1(n2834), .B2(n354), .A(n2392), .ZN(n2358) );
  AOI222_X2 U1374 ( .A1(n3142), .A2(n412), .B1(n325), .B2(n409), .C1(n380), 
        .C2(n406), .ZN(n2392) );
  XOR2_X2 U1375 ( .A(n2359), .B(n280), .Z(n1877) );
  OAI21_X4 U1376 ( .B1(n2835), .B2(n354), .A(n2393), .ZN(n2359) );
  AOI222_X2 U1377 ( .A1(n3143), .A2(n409), .B1(n325), .B2(n406), .C1(n380), 
        .C2(n403), .ZN(n2393) );
  XOR2_X2 U1378 ( .A(n2360), .B(n280), .Z(n1878) );
  OAI21_X4 U1379 ( .B1(n2836), .B2(n354), .A(n2394), .ZN(n2360) );
  AOI222_X2 U1380 ( .A1(n3143), .A2(n406), .B1(n325), .B2(n403), .C1(n380), 
        .C2(n400), .ZN(n2394) );
  XOR2_X2 U1381 ( .A(n2361), .B(n280), .Z(n1879) );
  OAI21_X4 U1382 ( .B1(n2837), .B2(n354), .A(n2395), .ZN(n2361) );
  AOI222_X2 U1383 ( .A1(n3142), .A2(n403), .B1(n325), .B2(n400), .C1(n380), 
        .C2(n397), .ZN(n2395) );
  XOR2_X2 U1384 ( .A(n2362), .B(n280), .Z(n1880) );
  OAI21_X4 U1385 ( .B1(n2838), .B2(n354), .A(n2396), .ZN(n2362) );
  AOI222_X2 U1386 ( .A1(n3143), .A2(n400), .B1(n325), .B2(n397), .C1(n380), 
        .C2(n393), .ZN(n2396) );
  XOR2_X2 U1387 ( .A(n2363), .B(n280), .Z(n1881) );
  OAI21_X4 U1388 ( .B1(n2839), .B2(n354), .A(n2397), .ZN(n2363) );
  AOI222_X2 U1389 ( .A1(n3142), .A2(n397), .B1(n325), .B2(n393), .C1(n380), 
        .C2(n390), .ZN(n2397) );
  XOR2_X2 U1390 ( .A(n2364), .B(n280), .Z(n1882) );
  OAI21_X4 U1391 ( .B1(n2840), .B2(n354), .A(n2398), .ZN(n2364) );
  OAI21_X4 U1394 ( .B1(n2841), .B2(n354), .A(n2399), .ZN(n2365) );
  AND2_X4 U1396 ( .A1(n3142), .A2(n390), .ZN(n1388) );
  XOR2_X2 U1398 ( .A(n2400), .B(n277), .Z(n1885) );
  OAI21_X4 U1399 ( .B1(n2808), .B2(n3126), .A(n2434), .ZN(n2400) );
  NAND2_X4 U1400 ( .A1(n378), .A2(n484), .ZN(n2434) );
  XOR2_X2 U1401 ( .A(n2401), .B(n277), .Z(n1886) );
  OAI21_X4 U1402 ( .B1(n2809), .B2(n3126), .A(n2435), .ZN(n2401) );
  AOI21_X4 U1403 ( .B1(n378), .B2(n481), .A(n1389), .ZN(n2435) );
  AND2_X4 U1404 ( .A1(n323), .A2(n484), .ZN(n1389) );
  XOR2_X2 U1405 ( .A(n2402), .B(n277), .Z(n1887) );
  OAI21_X4 U1406 ( .B1(n2810), .B2(n351), .A(n2436), .ZN(n2402) );
  AOI222_X2 U1407 ( .A1(n3146), .A2(n484), .B1(n323), .B2(n481), .C1(n378), 
        .C2(n478), .ZN(n2436) );
  XOR2_X2 U1408 ( .A(n2403), .B(n277), .Z(n1888) );
  OAI21_X4 U1409 ( .B1(n2811), .B2(n351), .A(n2437), .ZN(n2403) );
  AOI222_X2 U1410 ( .A1(n3145), .A2(n481), .B1(n323), .B2(n478), .C1(n378), 
        .C2(n475), .ZN(n2437) );
  XOR2_X2 U1411 ( .A(n2404), .B(n277), .Z(n1889) );
  OAI21_X4 U1412 ( .B1(n2812), .B2(n351), .A(n2438), .ZN(n2404) );
  AOI222_X2 U1413 ( .A1(n3146), .A2(n478), .B1(n323), .B2(n475), .C1(n378), 
        .C2(n472), .ZN(n2438) );
  XOR2_X2 U1414 ( .A(n2405), .B(n277), .Z(n1890) );
  OAI21_X4 U1415 ( .B1(n2813), .B2(n351), .A(n2439), .ZN(n2405) );
  AOI222_X2 U1416 ( .A1(n3145), .A2(n475), .B1(n323), .B2(n472), .C1(n378), 
        .C2(n469), .ZN(n2439) );
  XOR2_X2 U1417 ( .A(n2406), .B(n277), .Z(n1891) );
  OAI21_X4 U1418 ( .B1(n2814), .B2(n351), .A(n2440), .ZN(n2406) );
  AOI222_X2 U1419 ( .A1(n3146), .A2(n472), .B1(n323), .B2(n469), .C1(n378), 
        .C2(n466), .ZN(n2440) );
  XOR2_X2 U1420 ( .A(n2407), .B(n277), .Z(n1892) );
  OAI21_X4 U1421 ( .B1(n2815), .B2(n351), .A(n2441), .ZN(n2407) );
  AOI222_X2 U1422 ( .A1(n3145), .A2(n469), .B1(n323), .B2(n466), .C1(n378), 
        .C2(n463), .ZN(n2441) );
  XOR2_X2 U1423 ( .A(n2408), .B(n277), .Z(n1893) );
  OAI21_X4 U1424 ( .B1(n2816), .B2(n351), .A(n2442), .ZN(n2408) );
  AOI222_X2 U1425 ( .A1(n3146), .A2(n466), .B1(n323), .B2(n463), .C1(n378), 
        .C2(n460), .ZN(n2442) );
  XOR2_X2 U1426 ( .A(n2409), .B(n277), .Z(n1894) );
  OAI21_X4 U1427 ( .B1(n2817), .B2(n351), .A(n2443), .ZN(n2409) );
  AOI222_X2 U1428 ( .A1(n3145), .A2(n463), .B1(n323), .B2(n460), .C1(n378), 
        .C2(n457), .ZN(n2443) );
  XOR2_X2 U1429 ( .A(n2410), .B(n277), .Z(n1895) );
  OAI21_X4 U1430 ( .B1(n2818), .B2(n351), .A(n2444), .ZN(n2410) );
  AOI222_X2 U1431 ( .A1(n3146), .A2(n460), .B1(n323), .B2(n457), .C1(n378), 
        .C2(n454), .ZN(n2444) );
  XOR2_X2 U1432 ( .A(n2411), .B(n277), .Z(n1896) );
  OAI21_X4 U1433 ( .B1(n2819), .B2(n351), .A(n2445), .ZN(n2411) );
  AOI222_X2 U1434 ( .A1(n3145), .A2(n457), .B1(n323), .B2(n454), .C1(n378), 
        .C2(n451), .ZN(n2445) );
  XOR2_X2 U1435 ( .A(n2412), .B(n277), .Z(n1897) );
  OAI21_X4 U1436 ( .B1(n2820), .B2(n351), .A(n2446), .ZN(n2412) );
  AOI222_X2 U1437 ( .A1(n3145), .A2(n454), .B1(n323), .B2(n451), .C1(n378), 
        .C2(n448), .ZN(n2446) );
  XOR2_X2 U1438 ( .A(n2413), .B(n277), .Z(n1898) );
  OAI21_X4 U1439 ( .B1(n2821), .B2(n351), .A(n2447), .ZN(n2413) );
  AOI222_X2 U1440 ( .A1(n3146), .A2(n451), .B1(n323), .B2(n448), .C1(n378), 
        .C2(n445), .ZN(n2447) );
  XOR2_X2 U1441 ( .A(n2414), .B(n277), .Z(n1899) );
  OAI21_X4 U1442 ( .B1(n2822), .B2(n351), .A(n2448), .ZN(n2414) );
  AOI222_X2 U1443 ( .A1(n3146), .A2(n448), .B1(n323), .B2(n445), .C1(n378), 
        .C2(n442), .ZN(n2448) );
  XOR2_X2 U1444 ( .A(n2415), .B(n277), .Z(n1900) );
  OAI21_X4 U1445 ( .B1(n2823), .B2(n351), .A(n2449), .ZN(n2415) );
  AOI222_X2 U1446 ( .A1(n3146), .A2(n445), .B1(n323), .B2(n442), .C1(n378), 
        .C2(n439), .ZN(n2449) );
  XOR2_X2 U1447 ( .A(n2416), .B(n277), .Z(n1901) );
  OAI21_X4 U1448 ( .B1(n2824), .B2(n351), .A(n2450), .ZN(n2416) );
  AOI222_X2 U1449 ( .A1(n3145), .A2(n442), .B1(n323), .B2(n439), .C1(n378), 
        .C2(n436), .ZN(n2450) );
  XOR2_X2 U1450 ( .A(n2417), .B(n277), .Z(n1902) );
  OAI21_X4 U1451 ( .B1(n2825), .B2(n351), .A(n2451), .ZN(n2417) );
  AOI222_X2 U1452 ( .A1(n3145), .A2(n439), .B1(n323), .B2(n436), .C1(n378), 
        .C2(n433), .ZN(n2451) );
  XOR2_X2 U1453 ( .A(n2418), .B(n277), .Z(n1903) );
  OAI21_X4 U1454 ( .B1(n2826), .B2(n351), .A(n2452), .ZN(n2418) );
  AOI222_X2 U1455 ( .A1(n3145), .A2(n436), .B1(n323), .B2(n433), .C1(n378), 
        .C2(n430), .ZN(n2452) );
  XOR2_X2 U1456 ( .A(n2419), .B(n277), .Z(n1904) );
  OAI21_X4 U1457 ( .B1(n2827), .B2(n351), .A(n2453), .ZN(n2419) );
  AOI222_X2 U1458 ( .A1(n3146), .A2(n433), .B1(n323), .B2(n430), .C1(n378), 
        .C2(n427), .ZN(n2453) );
  XOR2_X2 U1459 ( .A(n2420), .B(n277), .Z(n1905) );
  OAI21_X4 U1460 ( .B1(n2828), .B2(n351), .A(n2454), .ZN(n2420) );
  AOI222_X2 U1461 ( .A1(n3146), .A2(n430), .B1(n323), .B2(n427), .C1(n378), 
        .C2(n424), .ZN(n2454) );
  XOR2_X2 U1462 ( .A(n2421), .B(n277), .Z(n1906) );
  OAI21_X4 U1463 ( .B1(n2829), .B2(n351), .A(n2455), .ZN(n2421) );
  AOI222_X2 U1464 ( .A1(n3145), .A2(n427), .B1(n323), .B2(n424), .C1(n378), 
        .C2(n421), .ZN(n2455) );
  XOR2_X2 U1465 ( .A(n2422), .B(n277), .Z(n1907) );
  OAI21_X4 U1466 ( .B1(n2830), .B2(n351), .A(n2456), .ZN(n2422) );
  AOI222_X2 U1467 ( .A1(n3145), .A2(n424), .B1(n323), .B2(n421), .C1(n378), 
        .C2(n418), .ZN(n2456) );
  XOR2_X2 U1468 ( .A(n2423), .B(n277), .Z(n1908) );
  OAI21_X4 U1469 ( .B1(n2831), .B2(n351), .A(n2457), .ZN(n2423) );
  AOI222_X2 U1470 ( .A1(n3146), .A2(n421), .B1(n323), .B2(n418), .C1(n378), 
        .C2(n415), .ZN(n2457) );
  XOR2_X2 U1471 ( .A(n2424), .B(n277), .Z(n1909) );
  OAI21_X4 U1472 ( .B1(n2832), .B2(n351), .A(n2458), .ZN(n2424) );
  AOI222_X2 U1473 ( .A1(n3145), .A2(n418), .B1(n323), .B2(n415), .C1(n378), 
        .C2(n412), .ZN(n2458) );
  XOR2_X2 U1474 ( .A(n2425), .B(n277), .Z(n1910) );
  OAI21_X4 U1475 ( .B1(n2833), .B2(n351), .A(n2459), .ZN(n2425) );
  AOI222_X2 U1476 ( .A1(n3146), .A2(n415), .B1(n323), .B2(n412), .C1(n378), 
        .C2(n409), .ZN(n2459) );
  XOR2_X2 U1477 ( .A(n2426), .B(n277), .Z(n1911) );
  OAI21_X4 U1478 ( .B1(n2834), .B2(n351), .A(n2460), .ZN(n2426) );
  AOI222_X2 U1479 ( .A1(n3146), .A2(n412), .B1(n323), .B2(n409), .C1(n378), 
        .C2(n406), .ZN(n2460) );
  XOR2_X2 U1480 ( .A(n2427), .B(n277), .Z(n1912) );
  OAI21_X4 U1481 ( .B1(n2835), .B2(n351), .A(n2461), .ZN(n2427) );
  AOI222_X2 U1482 ( .A1(n3145), .A2(n409), .B1(n323), .B2(n406), .C1(n378), 
        .C2(n403), .ZN(n2461) );
  XOR2_X2 U1483 ( .A(n2428), .B(n277), .Z(n1913) );
  OAI21_X4 U1484 ( .B1(n2836), .B2(n351), .A(n2462), .ZN(n2428) );
  AOI222_X2 U1485 ( .A1(n3146), .A2(n406), .B1(n323), .B2(n403), .C1(n378), 
        .C2(n400), .ZN(n2462) );
  XOR2_X2 U1486 ( .A(n2429), .B(n277), .Z(n1914) );
  OAI21_X4 U1487 ( .B1(n2837), .B2(n351), .A(n2463), .ZN(n2429) );
  AOI222_X2 U1488 ( .A1(n3145), .A2(n403), .B1(n323), .B2(n400), .C1(n378), 
        .C2(n397), .ZN(n2463) );
  XOR2_X2 U1489 ( .A(n2430), .B(n277), .Z(n1915) );
  OAI21_X4 U1490 ( .B1(n2838), .B2(n351), .A(n2464), .ZN(n2430) );
  AOI222_X2 U1491 ( .A1(n3146), .A2(n400), .B1(n323), .B2(n397), .C1(n378), 
        .C2(n393), .ZN(n2464) );
  XOR2_X2 U1492 ( .A(n2431), .B(n277), .Z(n1916) );
  OAI21_X4 U1493 ( .B1(n2839), .B2(n351), .A(n2465), .ZN(n2431) );
  AOI222_X2 U1494 ( .A1(n3145), .A2(n397), .B1(n323), .B2(n393), .C1(n378), 
        .C2(n390), .ZN(n2465) );
  XOR2_X2 U1495 ( .A(n2432), .B(n277), .Z(n1917) );
  OAI21_X4 U1496 ( .B1(n2840), .B2(n351), .A(n2466), .ZN(n2432) );
  XOR2_X2 U1498 ( .A(n2433), .B(n277), .Z(n1918) );
  OAI21_X4 U1499 ( .B1(n2841), .B2(n351), .A(n2467), .ZN(n2433) );
  AND2_X4 U1501 ( .A1(n3145), .A2(n390), .ZN(n1391) );
  XOR2_X2 U1503 ( .A(n2468), .B(n274), .Z(n1920) );
  OAI21_X4 U1504 ( .B1(n2808), .B2(n3127), .A(n2502), .ZN(n2468) );
  NAND2_X4 U1505 ( .A1(n376), .A2(n484), .ZN(n2502) );
  XOR2_X2 U1506 ( .A(n2469), .B(n274), .Z(n1921) );
  OAI21_X4 U1507 ( .B1(n2809), .B2(n3127), .A(n2503), .ZN(n2469) );
  AOI21_X4 U1508 ( .B1(n376), .B2(n481), .A(n1392), .ZN(n2503) );
  AND2_X4 U1509 ( .A1(n321), .A2(n484), .ZN(n1392) );
  XOR2_X2 U1510 ( .A(n2470), .B(n274), .Z(n1922) );
  OAI21_X4 U1511 ( .B1(n2810), .B2(n348), .A(n2504), .ZN(n2470) );
  AOI222_X2 U1512 ( .A1(n3149), .A2(n484), .B1(n321), .B2(n481), .C1(n376), 
        .C2(n478), .ZN(n2504) );
  XOR2_X2 U1513 ( .A(n2471), .B(n274), .Z(n1923) );
  OAI21_X4 U1514 ( .B1(n2811), .B2(n348), .A(n2505), .ZN(n2471) );
  AOI222_X2 U1515 ( .A1(n3148), .A2(n481), .B1(n321), .B2(n478), .C1(n376), 
        .C2(n475), .ZN(n2505) );
  XOR2_X2 U1516 ( .A(n2472), .B(n274), .Z(n1924) );
  OAI21_X4 U1517 ( .B1(n2812), .B2(n348), .A(n2506), .ZN(n2472) );
  AOI222_X2 U1518 ( .A1(n3149), .A2(n478), .B1(n321), .B2(n475), .C1(n376), 
        .C2(n472), .ZN(n2506) );
  XOR2_X2 U1519 ( .A(n2473), .B(n274), .Z(n1925) );
  OAI21_X4 U1520 ( .B1(n2813), .B2(n348), .A(n2507), .ZN(n2473) );
  AOI222_X2 U1521 ( .A1(n3148), .A2(n475), .B1(n321), .B2(n472), .C1(n376), 
        .C2(n469), .ZN(n2507) );
  XOR2_X2 U1522 ( .A(n2474), .B(n274), .Z(n1926) );
  OAI21_X4 U1523 ( .B1(n2814), .B2(n348), .A(n2508), .ZN(n2474) );
  AOI222_X2 U1524 ( .A1(n3149), .A2(n472), .B1(n321), .B2(n469), .C1(n376), 
        .C2(n466), .ZN(n2508) );
  XOR2_X2 U1525 ( .A(n2475), .B(n274), .Z(n1927) );
  OAI21_X4 U1526 ( .B1(n2815), .B2(n348), .A(n2509), .ZN(n2475) );
  AOI222_X2 U1527 ( .A1(n3148), .A2(n469), .B1(n321), .B2(n466), .C1(n376), 
        .C2(n463), .ZN(n2509) );
  XOR2_X2 U1528 ( .A(n2476), .B(n274), .Z(n1928) );
  OAI21_X4 U1529 ( .B1(n2816), .B2(n348), .A(n2510), .ZN(n2476) );
  AOI222_X2 U1530 ( .A1(n3149), .A2(n466), .B1(n321), .B2(n463), .C1(n376), 
        .C2(n460), .ZN(n2510) );
  XOR2_X2 U1531 ( .A(n2477), .B(n274), .Z(n1929) );
  OAI21_X4 U1532 ( .B1(n2817), .B2(n348), .A(n2511), .ZN(n2477) );
  AOI222_X2 U1533 ( .A1(n3148), .A2(n463), .B1(n321), .B2(n460), .C1(n376), 
        .C2(n457), .ZN(n2511) );
  XOR2_X2 U1534 ( .A(n2478), .B(n274), .Z(n1930) );
  OAI21_X4 U1535 ( .B1(n2818), .B2(n348), .A(n2512), .ZN(n2478) );
  AOI222_X2 U1536 ( .A1(n3148), .A2(n460), .B1(n321), .B2(n457), .C1(n376), 
        .C2(n454), .ZN(n2512) );
  XOR2_X2 U1537 ( .A(n2479), .B(n274), .Z(n1931) );
  OAI21_X4 U1538 ( .B1(n2819), .B2(n348), .A(n2513), .ZN(n2479) );
  AOI222_X2 U1539 ( .A1(n3149), .A2(n457), .B1(n321), .B2(n454), .C1(n376), 
        .C2(n451), .ZN(n2513) );
  XOR2_X2 U1540 ( .A(n2480), .B(n274), .Z(n1932) );
  OAI21_X4 U1541 ( .B1(n2820), .B2(n348), .A(n2514), .ZN(n2480) );
  AOI222_X2 U1542 ( .A1(n3149), .A2(n454), .B1(n321), .B2(n451), .C1(n376), 
        .C2(n448), .ZN(n2514) );
  XOR2_X2 U1543 ( .A(n2481), .B(n274), .Z(n1933) );
  OAI21_X4 U1544 ( .B1(n2821), .B2(n348), .A(n2515), .ZN(n2481) );
  AOI222_X2 U1545 ( .A1(n3148), .A2(n451), .B1(n321), .B2(n448), .C1(n376), 
        .C2(n445), .ZN(n2515) );
  XOR2_X2 U1546 ( .A(n2482), .B(n274), .Z(n1934) );
  OAI21_X4 U1547 ( .B1(n2822), .B2(n348), .A(n2516), .ZN(n2482) );
  AOI222_X2 U1548 ( .A1(n3149), .A2(n448), .B1(n321), .B2(n445), .C1(n376), 
        .C2(n442), .ZN(n2516) );
  XOR2_X2 U1549 ( .A(n2483), .B(n274), .Z(n1935) );
  OAI21_X4 U1550 ( .B1(n2823), .B2(n348), .A(n2517), .ZN(n2483) );
  AOI222_X2 U1551 ( .A1(n3148), .A2(n445), .B1(n321), .B2(n442), .C1(n376), 
        .C2(n439), .ZN(n2517) );
  XOR2_X2 U1552 ( .A(n2484), .B(n274), .Z(n1936) );
  OAI21_X4 U1553 ( .B1(n2824), .B2(n348), .A(n2518), .ZN(n2484) );
  AOI222_X2 U1554 ( .A1(n3149), .A2(n442), .B1(n321), .B2(n439), .C1(n376), 
        .C2(n436), .ZN(n2518) );
  XOR2_X2 U1555 ( .A(n2485), .B(n274), .Z(n1937) );
  OAI21_X4 U1556 ( .B1(n2825), .B2(n348), .A(n2519), .ZN(n2485) );
  AOI222_X2 U1557 ( .A1(n3149), .A2(n439), .B1(n321), .B2(n436), .C1(n376), 
        .C2(n433), .ZN(n2519) );
  XOR2_X2 U1558 ( .A(n2486), .B(n274), .Z(n1938) );
  OAI21_X4 U1559 ( .B1(n2826), .B2(n348), .A(n2520), .ZN(n2486) );
  AOI222_X2 U1560 ( .A1(n3148), .A2(n436), .B1(n321), .B2(n433), .C1(n376), 
        .C2(n430), .ZN(n2520) );
  XOR2_X2 U1561 ( .A(n2487), .B(n274), .Z(n1939) );
  OAI21_X4 U1562 ( .B1(n2827), .B2(n348), .A(n2521), .ZN(n2487) );
  AOI222_X2 U1563 ( .A1(n3149), .A2(n433), .B1(n321), .B2(n430), .C1(n376), 
        .C2(n427), .ZN(n2521) );
  XOR2_X2 U1564 ( .A(n2488), .B(n274), .Z(n1940) );
  OAI21_X4 U1565 ( .B1(n2828), .B2(n348), .A(n2522), .ZN(n2488) );
  AOI222_X2 U1566 ( .A1(n3148), .A2(n430), .B1(n321), .B2(n427), .C1(n376), 
        .C2(n424), .ZN(n2522) );
  XOR2_X2 U1567 ( .A(n2489), .B(n274), .Z(n1941) );
  OAI21_X4 U1568 ( .B1(n2829), .B2(n348), .A(n2523), .ZN(n2489) );
  AOI222_X2 U1569 ( .A1(n3149), .A2(n427), .B1(n321), .B2(n424), .C1(n376), 
        .C2(n421), .ZN(n2523) );
  XOR2_X2 U1570 ( .A(n2490), .B(n274), .Z(n1942) );
  OAI21_X4 U1571 ( .B1(n2830), .B2(n348), .A(n2524), .ZN(n2490) );
  AOI222_X2 U1572 ( .A1(n3148), .A2(n424), .B1(n321), .B2(n421), .C1(n376), 
        .C2(n418), .ZN(n2524) );
  XOR2_X2 U1573 ( .A(n2491), .B(n274), .Z(n1943) );
  OAI21_X4 U1574 ( .B1(n2831), .B2(n348), .A(n2525), .ZN(n2491) );
  AOI222_X2 U1575 ( .A1(n3149), .A2(n421), .B1(n321), .B2(n418), .C1(n376), 
        .C2(n415), .ZN(n2525) );
  XOR2_X2 U1576 ( .A(n2492), .B(n274), .Z(n1944) );
  OAI21_X4 U1577 ( .B1(n2832), .B2(n348), .A(n2526), .ZN(n2492) );
  AOI222_X2 U1578 ( .A1(n3148), .A2(n418), .B1(n321), .B2(n415), .C1(n376), 
        .C2(n412), .ZN(n2526) );
  XOR2_X2 U1579 ( .A(n2493), .B(n274), .Z(n1945) );
  OAI21_X4 U1580 ( .B1(n2833), .B2(n348), .A(n2527), .ZN(n2493) );
  AOI222_X2 U1581 ( .A1(n3148), .A2(n415), .B1(n321), .B2(n412), .C1(n376), 
        .C2(n409), .ZN(n2527) );
  XOR2_X2 U1582 ( .A(n2494), .B(n274), .Z(n1946) );
  OAI21_X4 U1583 ( .B1(n2834), .B2(n348), .A(n2528), .ZN(n2494) );
  AOI222_X2 U1584 ( .A1(n3149), .A2(n412), .B1(n321), .B2(n409), .C1(n376), 
        .C2(n406), .ZN(n2528) );
  XOR2_X2 U1585 ( .A(n2495), .B(n274), .Z(n1947) );
  OAI21_X4 U1586 ( .B1(n2835), .B2(n348), .A(n2529), .ZN(n2495) );
  AOI222_X2 U1587 ( .A1(n3148), .A2(n409), .B1(n321), .B2(n406), .C1(n376), 
        .C2(n403), .ZN(n2529) );
  XOR2_X2 U1588 ( .A(n2496), .B(n274), .Z(n1948) );
  OAI21_X4 U1589 ( .B1(n2836), .B2(n348), .A(n2530), .ZN(n2496) );
  AOI222_X2 U1590 ( .A1(n3149), .A2(n406), .B1(n321), .B2(n403), .C1(n376), 
        .C2(n400), .ZN(n2530) );
  XOR2_X2 U1591 ( .A(n2497), .B(n274), .Z(n1949) );
  OAI21_X4 U1592 ( .B1(n2837), .B2(n348), .A(n2531), .ZN(n2497) );
  AOI222_X2 U1593 ( .A1(n3148), .A2(n403), .B1(n321), .B2(n400), .C1(n376), 
        .C2(n397), .ZN(n2531) );
  XOR2_X2 U1594 ( .A(n2498), .B(n274), .Z(n1950) );
  OAI21_X4 U1595 ( .B1(n2838), .B2(n348), .A(n2532), .ZN(n2498) );
  AOI222_X2 U1596 ( .A1(n3149), .A2(n400), .B1(n321), .B2(n397), .C1(n376), 
        .C2(n393), .ZN(n2532) );
  XOR2_X2 U1597 ( .A(n2499), .B(n274), .Z(n1951) );
  OAI21_X4 U1598 ( .B1(n2839), .B2(n348), .A(n2533), .ZN(n2499) );
  AOI222_X2 U1599 ( .A1(n3148), .A2(n397), .B1(n321), .B2(n393), .C1(n376), 
        .C2(n390), .ZN(n2533) );
  XOR2_X2 U1600 ( .A(n2500), .B(n274), .Z(n1952) );
  OAI21_X4 U1601 ( .B1(n2840), .B2(n348), .A(n2534), .ZN(n2500) );
  XOR2_X2 U1603 ( .A(n2501), .B(n274), .Z(n1953) );
  OAI21_X4 U1604 ( .B1(n2841), .B2(n348), .A(n2535), .ZN(n2501) );
  AND2_X4 U1606 ( .A1(n3148), .A2(n390), .ZN(n1394) );
  XOR2_X2 U1608 ( .A(n2536), .B(n271), .Z(n1955) );
  OAI21_X4 U1609 ( .B1(n2808), .B2(n345), .A(n2570), .ZN(n2536) );
  NAND2_X4 U1610 ( .A1(n374), .A2(n484), .ZN(n2570) );
  XOR2_X2 U1611 ( .A(n2537), .B(n271), .Z(n1956) );
  OAI21_X4 U1612 ( .B1(n2809), .B2(n345), .A(n2571), .ZN(n2537) );
  AOI21_X4 U1613 ( .B1(n374), .B2(n481), .A(n1395), .ZN(n2571) );
  AND2_X4 U1614 ( .A1(n319), .A2(n484), .ZN(n1395) );
  XOR2_X2 U1615 ( .A(n2538), .B(n271), .Z(n1957) );
  OAI21_X4 U1616 ( .B1(n2810), .B2(n345), .A(n2572), .ZN(n2538) );
  AOI222_X2 U1617 ( .A1(n297), .A2(n484), .B1(n319), .B2(n481), .C1(n374), 
        .C2(n478), .ZN(n2572) );
  XOR2_X2 U1618 ( .A(n2539), .B(n271), .Z(n1958) );
  OAI21_X4 U1619 ( .B1(n2811), .B2(n345), .A(n2573), .ZN(n2539) );
  AOI222_X2 U1620 ( .A1(n297), .A2(n481), .B1(n319), .B2(n478), .C1(n374), 
        .C2(n475), .ZN(n2573) );
  XOR2_X2 U1621 ( .A(n2540), .B(n271), .Z(n1959) );
  OAI21_X4 U1622 ( .B1(n2812), .B2(n345), .A(n2574), .ZN(n2540) );
  AOI222_X2 U1623 ( .A1(n297), .A2(n478), .B1(n319), .B2(n475), .C1(n374), 
        .C2(n472), .ZN(n2574) );
  XOR2_X2 U1624 ( .A(n2541), .B(n271), .Z(n1960) );
  OAI21_X4 U1625 ( .B1(n2813), .B2(n345), .A(n2575), .ZN(n2541) );
  AOI222_X2 U1626 ( .A1(n297), .A2(n475), .B1(n319), .B2(n472), .C1(n374), 
        .C2(n469), .ZN(n2575) );
  XOR2_X2 U1627 ( .A(n2542), .B(n271), .Z(n1961) );
  OAI21_X4 U1628 ( .B1(n2814), .B2(n345), .A(n2576), .ZN(n2542) );
  AOI222_X2 U1629 ( .A1(n297), .A2(n472), .B1(n319), .B2(n469), .C1(n374), 
        .C2(n466), .ZN(n2576) );
  XOR2_X2 U1630 ( .A(n2543), .B(n271), .Z(n1962) );
  OAI21_X4 U1631 ( .B1(n2815), .B2(n345), .A(n2577), .ZN(n2543) );
  AOI222_X2 U1632 ( .A1(n297), .A2(n469), .B1(n319), .B2(n466), .C1(n374), 
        .C2(n463), .ZN(n2577) );
  XOR2_X2 U1633 ( .A(n2544), .B(n271), .Z(n1963) );
  OAI21_X4 U1634 ( .B1(n2816), .B2(n345), .A(n2578), .ZN(n2544) );
  AOI222_X2 U1635 ( .A1(n297), .A2(n466), .B1(n319), .B2(n463), .C1(n374), 
        .C2(n460), .ZN(n2578) );
  XOR2_X2 U1636 ( .A(n2545), .B(n271), .Z(n1964) );
  OAI21_X4 U1637 ( .B1(n2817), .B2(n345), .A(n2579), .ZN(n2545) );
  AOI222_X2 U1638 ( .A1(n297), .A2(n463), .B1(n319), .B2(n460), .C1(n374), 
        .C2(n457), .ZN(n2579) );
  XOR2_X2 U1639 ( .A(n2546), .B(n271), .Z(n1965) );
  OAI21_X4 U1640 ( .B1(n2818), .B2(n345), .A(n2580), .ZN(n2546) );
  AOI222_X2 U1641 ( .A1(n297), .A2(n460), .B1(n319), .B2(n457), .C1(n374), 
        .C2(n454), .ZN(n2580) );
  XOR2_X2 U1642 ( .A(n2547), .B(n271), .Z(n1966) );
  OAI21_X4 U1643 ( .B1(n2819), .B2(n345), .A(n2581), .ZN(n2547) );
  AOI222_X2 U1644 ( .A1(n297), .A2(n457), .B1(n319), .B2(n454), .C1(n374), 
        .C2(n451), .ZN(n2581) );
  XOR2_X2 U1645 ( .A(n2548), .B(n271), .Z(n1967) );
  OAI21_X4 U1646 ( .B1(n2820), .B2(n345), .A(n2582), .ZN(n2548) );
  AOI222_X2 U1647 ( .A1(n297), .A2(n454), .B1(n319), .B2(n451), .C1(n374), 
        .C2(n448), .ZN(n2582) );
  XOR2_X2 U1648 ( .A(n2549), .B(n271), .Z(n1968) );
  OAI21_X4 U1649 ( .B1(n2821), .B2(n345), .A(n2583), .ZN(n2549) );
  AOI222_X2 U1650 ( .A1(n297), .A2(n451), .B1(n319), .B2(n448), .C1(n374), 
        .C2(n445), .ZN(n2583) );
  XOR2_X2 U1651 ( .A(n2550), .B(n271), .Z(n1969) );
  OAI21_X4 U1652 ( .B1(n2822), .B2(n345), .A(n2584), .ZN(n2550) );
  AOI222_X2 U1653 ( .A1(n297), .A2(n448), .B1(n319), .B2(n445), .C1(n374), 
        .C2(n442), .ZN(n2584) );
  XOR2_X2 U1654 ( .A(n2551), .B(n271), .Z(n1970) );
  OAI21_X4 U1655 ( .B1(n2823), .B2(n345), .A(n2585), .ZN(n2551) );
  AOI222_X2 U1656 ( .A1(n297), .A2(n445), .B1(n319), .B2(n442), .C1(n374), 
        .C2(n439), .ZN(n2585) );
  XOR2_X2 U1657 ( .A(n2552), .B(n271), .Z(n1971) );
  OAI21_X4 U1658 ( .B1(n2824), .B2(n345), .A(n2586), .ZN(n2552) );
  AOI222_X2 U1659 ( .A1(n297), .A2(n442), .B1(n319), .B2(n439), .C1(n374), 
        .C2(n436), .ZN(n2586) );
  XOR2_X2 U1660 ( .A(n2553), .B(n271), .Z(n1972) );
  OAI21_X4 U1661 ( .B1(n2825), .B2(n345), .A(n2587), .ZN(n2553) );
  AOI222_X2 U1662 ( .A1(n297), .A2(n439), .B1(n319), .B2(n436), .C1(n374), 
        .C2(n433), .ZN(n2587) );
  XOR2_X2 U1663 ( .A(n2554), .B(n271), .Z(n1973) );
  OAI21_X4 U1664 ( .B1(n2826), .B2(n345), .A(n2588), .ZN(n2554) );
  AOI222_X2 U1665 ( .A1(n297), .A2(n436), .B1(n319), .B2(n433), .C1(n374), 
        .C2(n430), .ZN(n2588) );
  XOR2_X2 U1666 ( .A(n2555), .B(n271), .Z(n1974) );
  OAI21_X4 U1667 ( .B1(n2827), .B2(n345), .A(n2589), .ZN(n2555) );
  AOI222_X2 U1668 ( .A1(n297), .A2(n433), .B1(n319), .B2(n430), .C1(n374), 
        .C2(n427), .ZN(n2589) );
  XOR2_X2 U1669 ( .A(n2556), .B(n271), .Z(n1975) );
  OAI21_X4 U1670 ( .B1(n2828), .B2(n345), .A(n2590), .ZN(n2556) );
  AOI222_X2 U1671 ( .A1(n297), .A2(n430), .B1(n319), .B2(n427), .C1(n374), 
        .C2(n424), .ZN(n2590) );
  XOR2_X2 U1672 ( .A(n2557), .B(n271), .Z(n1976) );
  OAI21_X4 U1673 ( .B1(n2829), .B2(n345), .A(n2591), .ZN(n2557) );
  AOI222_X2 U1674 ( .A1(n297), .A2(n427), .B1(n319), .B2(n424), .C1(n374), 
        .C2(n421), .ZN(n2591) );
  XOR2_X2 U1675 ( .A(n2558), .B(n271), .Z(n1977) );
  OAI21_X4 U1676 ( .B1(n2830), .B2(n345), .A(n2592), .ZN(n2558) );
  AOI222_X2 U1677 ( .A1(n297), .A2(n424), .B1(n319), .B2(n421), .C1(n374), 
        .C2(n418), .ZN(n2592) );
  XOR2_X2 U1678 ( .A(n2559), .B(n271), .Z(n1978) );
  OAI21_X4 U1679 ( .B1(n2831), .B2(n345), .A(n2593), .ZN(n2559) );
  AOI222_X2 U1680 ( .A1(n297), .A2(n421), .B1(n319), .B2(n418), .C1(n374), 
        .C2(n415), .ZN(n2593) );
  XOR2_X2 U1681 ( .A(n2560), .B(n271), .Z(n1979) );
  OAI21_X4 U1682 ( .B1(n2832), .B2(n345), .A(n2594), .ZN(n2560) );
  AOI222_X2 U1683 ( .A1(n297), .A2(n418), .B1(n319), .B2(n415), .C1(n374), 
        .C2(n412), .ZN(n2594) );
  XOR2_X2 U1684 ( .A(n2561), .B(n271), .Z(n1980) );
  OAI21_X4 U1685 ( .B1(n2833), .B2(n345), .A(n2595), .ZN(n2561) );
  AOI222_X2 U1686 ( .A1(n297), .A2(n415), .B1(n319), .B2(n412), .C1(n374), 
        .C2(n409), .ZN(n2595) );
  XOR2_X2 U1687 ( .A(n2562), .B(n271), .Z(n1981) );
  OAI21_X4 U1688 ( .B1(n2834), .B2(n345), .A(n2596), .ZN(n2562) );
  AOI222_X2 U1689 ( .A1(n297), .A2(n412), .B1(n319), .B2(n409), .C1(n374), 
        .C2(n406), .ZN(n2596) );
  XOR2_X2 U1690 ( .A(n2563), .B(n271), .Z(n1982) );
  OAI21_X4 U1691 ( .B1(n2835), .B2(n345), .A(n2597), .ZN(n2563) );
  AOI222_X2 U1692 ( .A1(n297), .A2(n409), .B1(n319), .B2(n406), .C1(n374), 
        .C2(n403), .ZN(n2597) );
  XOR2_X2 U1693 ( .A(n2564), .B(n271), .Z(n1983) );
  OAI21_X4 U1694 ( .B1(n2836), .B2(n345), .A(n2598), .ZN(n2564) );
  AOI222_X2 U1695 ( .A1(n297), .A2(n406), .B1(n319), .B2(n403), .C1(n374), 
        .C2(n400), .ZN(n2598) );
  XOR2_X2 U1696 ( .A(n2565), .B(n271), .Z(n1984) );
  OAI21_X4 U1697 ( .B1(n2837), .B2(n345), .A(n2599), .ZN(n2565) );
  AOI222_X2 U1698 ( .A1(n297), .A2(n403), .B1(n319), .B2(n400), .C1(n374), 
        .C2(n397), .ZN(n2599) );
  XOR2_X2 U1699 ( .A(n2566), .B(n271), .Z(n1985) );
  OAI21_X4 U1700 ( .B1(n2838), .B2(n345), .A(n2600), .ZN(n2566) );
  AOI222_X2 U1701 ( .A1(n297), .A2(n400), .B1(n319), .B2(n397), .C1(n374), 
        .C2(n393), .ZN(n2600) );
  XOR2_X2 U1702 ( .A(n2567), .B(n271), .Z(n1986) );
  OAI21_X4 U1703 ( .B1(n2839), .B2(n345), .A(n2601), .ZN(n2567) );
  AOI222_X2 U1704 ( .A1(n297), .A2(n397), .B1(n319), .B2(n393), .C1(n374), 
        .C2(n390), .ZN(n2601) );
  XOR2_X2 U1705 ( .A(n2568), .B(n271), .Z(n1987) );
  OAI21_X4 U1706 ( .B1(n2840), .B2(n345), .A(n2602), .ZN(n2568) );
  AND2_X4 U1711 ( .A1(n297), .A2(n390), .ZN(n1397) );
  XOR2_X2 U1713 ( .A(n2604), .B(n268), .Z(n1990) );
  OAI21_X4 U1714 ( .B1(n2808), .B2(n342), .A(n2638), .ZN(n2604) );
  NAND2_X4 U1715 ( .A1(n372), .A2(n484), .ZN(n2638) );
  XOR2_X2 U1716 ( .A(n2605), .B(n268), .Z(n1991) );
  OAI21_X4 U1717 ( .B1(n2809), .B2(n342), .A(n2639), .ZN(n2605) );
  AOI21_X4 U1718 ( .B1(n372), .B2(n481), .A(n1398), .ZN(n2639) );
  AND2_X4 U1719 ( .A1(n317), .A2(n484), .ZN(n1398) );
  XOR2_X2 U1720 ( .A(n2606), .B(n268), .Z(n1992) );
  OAI21_X4 U1721 ( .B1(n2810), .B2(n342), .A(n2640), .ZN(n2606) );
  AOI222_X2 U1722 ( .A1(n295), .A2(n484), .B1(n317), .B2(n481), .C1(n372), 
        .C2(n478), .ZN(n2640) );
  XOR2_X2 U1723 ( .A(n2607), .B(n268), .Z(n1993) );
  OAI21_X4 U1724 ( .B1(n2811), .B2(n342), .A(n2641), .ZN(n2607) );
  AOI222_X2 U1725 ( .A1(n295), .A2(n481), .B1(n317), .B2(n478), .C1(n372), 
        .C2(n475), .ZN(n2641) );
  XOR2_X2 U1726 ( .A(n2608), .B(n268), .Z(n1994) );
  OAI21_X4 U1727 ( .B1(n2812), .B2(n342), .A(n2642), .ZN(n2608) );
  AOI222_X2 U1728 ( .A1(n295), .A2(n478), .B1(n317), .B2(n475), .C1(n372), 
        .C2(n472), .ZN(n2642) );
  XOR2_X2 U1729 ( .A(n2609), .B(n268), .Z(n1995) );
  OAI21_X4 U1730 ( .B1(n2813), .B2(n342), .A(n2643), .ZN(n2609) );
  AOI222_X2 U1731 ( .A1(n295), .A2(n475), .B1(n317), .B2(n472), .C1(n372), 
        .C2(n469), .ZN(n2643) );
  XOR2_X2 U1732 ( .A(n2610), .B(n268), .Z(n1996) );
  OAI21_X4 U1733 ( .B1(n2814), .B2(n342), .A(n2644), .ZN(n2610) );
  AOI222_X2 U1734 ( .A1(n295), .A2(n472), .B1(n317), .B2(n469), .C1(n372), 
        .C2(n466), .ZN(n2644) );
  XOR2_X2 U1735 ( .A(n2611), .B(n268), .Z(n1997) );
  OAI21_X4 U1736 ( .B1(n2815), .B2(n342), .A(n2645), .ZN(n2611) );
  AOI222_X2 U1737 ( .A1(n295), .A2(n469), .B1(n317), .B2(n466), .C1(n372), 
        .C2(n463), .ZN(n2645) );
  XOR2_X2 U1738 ( .A(n2612), .B(n268), .Z(n1998) );
  OAI21_X4 U1739 ( .B1(n2816), .B2(n342), .A(n2646), .ZN(n2612) );
  AOI222_X2 U1740 ( .A1(n295), .A2(n466), .B1(n317), .B2(n463), .C1(n372), 
        .C2(n460), .ZN(n2646) );
  XOR2_X2 U1741 ( .A(n2613), .B(n268), .Z(n1999) );
  OAI21_X4 U1742 ( .B1(n2817), .B2(n342), .A(n2647), .ZN(n2613) );
  AOI222_X2 U1743 ( .A1(n295), .A2(n463), .B1(n317), .B2(n460), .C1(n372), 
        .C2(n457), .ZN(n2647) );
  XOR2_X2 U1744 ( .A(n2614), .B(n268), .Z(n2000) );
  OAI21_X4 U1745 ( .B1(n2818), .B2(n342), .A(n2648), .ZN(n2614) );
  AOI222_X2 U1746 ( .A1(n295), .A2(n460), .B1(n317), .B2(n457), .C1(n372), 
        .C2(n454), .ZN(n2648) );
  XOR2_X2 U1747 ( .A(n2615), .B(n268), .Z(n2001) );
  OAI21_X4 U1748 ( .B1(n2819), .B2(n342), .A(n2649), .ZN(n2615) );
  AOI222_X2 U1749 ( .A1(n295), .A2(n457), .B1(n317), .B2(n454), .C1(n372), 
        .C2(n451), .ZN(n2649) );
  XOR2_X2 U1750 ( .A(n2616), .B(n268), .Z(n2002) );
  OAI21_X4 U1751 ( .B1(n2820), .B2(n342), .A(n2650), .ZN(n2616) );
  AOI222_X2 U1752 ( .A1(n295), .A2(n454), .B1(n317), .B2(n451), .C1(n372), 
        .C2(n448), .ZN(n2650) );
  XOR2_X2 U1753 ( .A(n2617), .B(n268), .Z(n2003) );
  OAI21_X4 U1754 ( .B1(n2821), .B2(n342), .A(n2651), .ZN(n2617) );
  AOI222_X2 U1755 ( .A1(n295), .A2(n451), .B1(n317), .B2(n448), .C1(n372), 
        .C2(n445), .ZN(n2651) );
  XOR2_X2 U1756 ( .A(n2618), .B(n268), .Z(n2004) );
  OAI21_X4 U1757 ( .B1(n2822), .B2(n342), .A(n2652), .ZN(n2618) );
  AOI222_X2 U1758 ( .A1(n295), .A2(n448), .B1(n317), .B2(n445), .C1(n372), 
        .C2(n442), .ZN(n2652) );
  XOR2_X2 U1759 ( .A(n2619), .B(n268), .Z(n2005) );
  OAI21_X4 U1760 ( .B1(n2823), .B2(n342), .A(n2653), .ZN(n2619) );
  AOI222_X2 U1761 ( .A1(n295), .A2(n445), .B1(n317), .B2(n442), .C1(n372), 
        .C2(n439), .ZN(n2653) );
  XOR2_X2 U1762 ( .A(n2620), .B(n268), .Z(n2006) );
  OAI21_X4 U1763 ( .B1(n2824), .B2(n342), .A(n2654), .ZN(n2620) );
  AOI222_X2 U1764 ( .A1(n295), .A2(n442), .B1(n317), .B2(n439), .C1(n372), 
        .C2(n436), .ZN(n2654) );
  XOR2_X2 U1765 ( .A(n2621), .B(n268), .Z(n2007) );
  OAI21_X4 U1766 ( .B1(n2825), .B2(n342), .A(n2655), .ZN(n2621) );
  AOI222_X2 U1767 ( .A1(n295), .A2(n439), .B1(n317), .B2(n436), .C1(n372), 
        .C2(n433), .ZN(n2655) );
  XOR2_X2 U1768 ( .A(n2622), .B(n268), .Z(n2008) );
  OAI21_X4 U1769 ( .B1(n2826), .B2(n342), .A(n2656), .ZN(n2622) );
  AOI222_X2 U1770 ( .A1(n295), .A2(n436), .B1(n317), .B2(n433), .C1(n372), 
        .C2(n430), .ZN(n2656) );
  XOR2_X2 U1771 ( .A(n2623), .B(n268), .Z(n2009) );
  OAI21_X4 U1772 ( .B1(n2827), .B2(n342), .A(n2657), .ZN(n2623) );
  AOI222_X2 U1773 ( .A1(n295), .A2(n433), .B1(n317), .B2(n430), .C1(n372), 
        .C2(n427), .ZN(n2657) );
  XOR2_X2 U1774 ( .A(n2624), .B(n268), .Z(n2010) );
  OAI21_X4 U1775 ( .B1(n2828), .B2(n342), .A(n2658), .ZN(n2624) );
  AOI222_X2 U1776 ( .A1(n295), .A2(n430), .B1(n317), .B2(n427), .C1(n372), 
        .C2(n424), .ZN(n2658) );
  XOR2_X2 U1777 ( .A(n2625), .B(n268), .Z(n2011) );
  OAI21_X4 U1778 ( .B1(n2829), .B2(n342), .A(n2659), .ZN(n2625) );
  AOI222_X2 U1779 ( .A1(n295), .A2(n427), .B1(n317), .B2(n424), .C1(n372), 
        .C2(n421), .ZN(n2659) );
  XOR2_X2 U1780 ( .A(n2626), .B(n268), .Z(n2012) );
  OAI21_X4 U1781 ( .B1(n2830), .B2(n342), .A(n2660), .ZN(n2626) );
  AOI222_X2 U1782 ( .A1(n295), .A2(n424), .B1(n317), .B2(n421), .C1(n372), 
        .C2(n418), .ZN(n2660) );
  XOR2_X2 U1783 ( .A(n2627), .B(n268), .Z(n2013) );
  OAI21_X4 U1784 ( .B1(n2831), .B2(n342), .A(n2661), .ZN(n2627) );
  AOI222_X2 U1785 ( .A1(n295), .A2(n421), .B1(n317), .B2(n418), .C1(n372), 
        .C2(n415), .ZN(n2661) );
  XOR2_X2 U1786 ( .A(n2628), .B(n268), .Z(n2014) );
  OAI21_X4 U1787 ( .B1(n2832), .B2(n342), .A(n2662), .ZN(n2628) );
  AOI222_X2 U1788 ( .A1(n295), .A2(n418), .B1(n317), .B2(n415), .C1(n372), 
        .C2(n412), .ZN(n2662) );
  XOR2_X2 U1789 ( .A(n2629), .B(n268), .Z(n2015) );
  OAI21_X4 U1790 ( .B1(n2833), .B2(n342), .A(n2663), .ZN(n2629) );
  AOI222_X2 U1791 ( .A1(n295), .A2(n415), .B1(n317), .B2(n412), .C1(n372), 
        .C2(n409), .ZN(n2663) );
  XOR2_X2 U1792 ( .A(n2630), .B(n268), .Z(n2016) );
  OAI21_X4 U1793 ( .B1(n2834), .B2(n342), .A(n2664), .ZN(n2630) );
  AOI222_X2 U1794 ( .A1(n295), .A2(n412), .B1(n317), .B2(n409), .C1(n372), 
        .C2(n406), .ZN(n2664) );
  XOR2_X2 U1795 ( .A(n2631), .B(n268), .Z(n2017) );
  OAI21_X4 U1796 ( .B1(n2835), .B2(n342), .A(n2665), .ZN(n2631) );
  AOI222_X2 U1797 ( .A1(n295), .A2(n409), .B1(n317), .B2(n406), .C1(n372), 
        .C2(n403), .ZN(n2665) );
  XOR2_X2 U1798 ( .A(n2632), .B(n268), .Z(n2018) );
  OAI21_X4 U1799 ( .B1(n2836), .B2(n342), .A(n2666), .ZN(n2632) );
  AOI222_X2 U1800 ( .A1(n295), .A2(n406), .B1(n317), .B2(n403), .C1(n372), 
        .C2(n400), .ZN(n2666) );
  XOR2_X2 U1801 ( .A(n2633), .B(n268), .Z(n2019) );
  OAI21_X4 U1802 ( .B1(n2837), .B2(n342), .A(n2667), .ZN(n2633) );
  AOI222_X2 U1803 ( .A1(n295), .A2(n403), .B1(n317), .B2(n400), .C1(n372), 
        .C2(n397), .ZN(n2667) );
  XOR2_X2 U1804 ( .A(n2634), .B(n268), .Z(n2020) );
  OAI21_X4 U1805 ( .B1(n2838), .B2(n342), .A(n2668), .ZN(n2634) );
  AOI222_X2 U1806 ( .A1(n295), .A2(n400), .B1(n317), .B2(n397), .C1(n372), 
        .C2(n393), .ZN(n2668) );
  XOR2_X2 U1807 ( .A(n2635), .B(n268), .Z(n2021) );
  OAI21_X4 U1808 ( .B1(n2839), .B2(n342), .A(n2669), .ZN(n2635) );
  AOI222_X2 U1809 ( .A1(n295), .A2(n397), .B1(n317), .B2(n393), .C1(n372), 
        .C2(n390), .ZN(n2669) );
  AND2_X4 U1816 ( .A1(n295), .A2(n390), .ZN(n1400) );
  XOR2_X2 U1818 ( .A(n2672), .B(n265), .Z(n2025) );
  OAI21_X4 U1819 ( .B1(n2808), .B2(n339), .A(n2706), .ZN(n2672) );
  NAND2_X4 U1820 ( .A1(n370), .A2(n484), .ZN(n2706) );
  XOR2_X2 U1821 ( .A(n2673), .B(n265), .Z(n2026) );
  OAI21_X4 U1822 ( .B1(n2809), .B2(n339), .A(n2707), .ZN(n2673) );
  AOI21_X4 U1823 ( .B1(n370), .B2(n481), .A(n1401), .ZN(n2707) );
  AND2_X4 U1824 ( .A1(n315), .A2(n484), .ZN(n1401) );
  XOR2_X2 U1825 ( .A(n2674), .B(n265), .Z(n2027) );
  OAI21_X4 U1826 ( .B1(n2810), .B2(n339), .A(n2708), .ZN(n2674) );
  AOI222_X2 U1827 ( .A1(n3217), .A2(n484), .B1(n315), .B2(n481), .C1(n370), 
        .C2(n478), .ZN(n2708) );
  XOR2_X2 U1828 ( .A(n2675), .B(n265), .Z(n2028) );
  OAI21_X4 U1829 ( .B1(n2811), .B2(n339), .A(n2709), .ZN(n2675) );
  AOI222_X2 U1830 ( .A1(n3217), .A2(n481), .B1(n315), .B2(n478), .C1(n370), 
        .C2(n475), .ZN(n2709) );
  XOR2_X2 U1831 ( .A(n2676), .B(n265), .Z(n2029) );
  OAI21_X4 U1832 ( .B1(n2812), .B2(n339), .A(n2710), .ZN(n2676) );
  AOI222_X2 U1833 ( .A1(n3217), .A2(n478), .B1(n315), .B2(n475), .C1(n370), 
        .C2(n472), .ZN(n2710) );
  XOR2_X2 U1834 ( .A(n2677), .B(n265), .Z(n2030) );
  OAI21_X4 U1835 ( .B1(n2813), .B2(n339), .A(n2711), .ZN(n2677) );
  AOI222_X2 U1836 ( .A1(n3217), .A2(n475), .B1(n315), .B2(n472), .C1(n370), 
        .C2(n469), .ZN(n2711) );
  XOR2_X2 U1837 ( .A(n2678), .B(n265), .Z(n2031) );
  OAI21_X4 U1838 ( .B1(n2814), .B2(n339), .A(n2712), .ZN(n2678) );
  AOI222_X2 U1839 ( .A1(n3217), .A2(n472), .B1(n315), .B2(n469), .C1(n370), 
        .C2(n466), .ZN(n2712) );
  XOR2_X2 U1840 ( .A(n2679), .B(n265), .Z(n2032) );
  OAI21_X4 U1841 ( .B1(n2815), .B2(n339), .A(n2713), .ZN(n2679) );
  AOI222_X2 U1842 ( .A1(n3217), .A2(n469), .B1(n315), .B2(n466), .C1(n370), 
        .C2(n463), .ZN(n2713) );
  XOR2_X2 U1843 ( .A(n2680), .B(n265), .Z(n2033) );
  OAI21_X4 U1844 ( .B1(n2816), .B2(n339), .A(n2714), .ZN(n2680) );
  AOI222_X2 U1845 ( .A1(n3217), .A2(n466), .B1(n315), .B2(n463), .C1(n370), 
        .C2(n460), .ZN(n2714) );
  XOR2_X2 U1846 ( .A(n2681), .B(n265), .Z(n2034) );
  OAI21_X4 U1847 ( .B1(n2817), .B2(n339), .A(n2715), .ZN(n2681) );
  AOI222_X2 U1848 ( .A1(n3217), .A2(n463), .B1(n315), .B2(n460), .C1(n370), 
        .C2(n457), .ZN(n2715) );
  XOR2_X2 U1849 ( .A(n2682), .B(n265), .Z(n2035) );
  OAI21_X4 U1850 ( .B1(n2818), .B2(n339), .A(n2716), .ZN(n2682) );
  AOI222_X2 U1851 ( .A1(n3217), .A2(n460), .B1(n315), .B2(n457), .C1(n370), 
        .C2(n454), .ZN(n2716) );
  XOR2_X2 U1852 ( .A(n2683), .B(n265), .Z(n2036) );
  OAI21_X4 U1853 ( .B1(n2819), .B2(n339), .A(n2717), .ZN(n2683) );
  AOI222_X2 U1854 ( .A1(n3217), .A2(n457), .B1(n315), .B2(n454), .C1(n370), 
        .C2(n451), .ZN(n2717) );
  XOR2_X2 U1855 ( .A(n2684), .B(n265), .Z(n2037) );
  OAI21_X4 U1856 ( .B1(n2820), .B2(n339), .A(n2718), .ZN(n2684) );
  AOI222_X2 U1857 ( .A1(n3217), .A2(n454), .B1(n315), .B2(n451), .C1(n370), 
        .C2(n448), .ZN(n2718) );
  XOR2_X2 U1858 ( .A(n2685), .B(n265), .Z(n2038) );
  OAI21_X4 U1859 ( .B1(n2821), .B2(n339), .A(n2719), .ZN(n2685) );
  AOI222_X2 U1860 ( .A1(n3217), .A2(n451), .B1(n315), .B2(n448), .C1(n370), 
        .C2(n445), .ZN(n2719) );
  XOR2_X2 U1861 ( .A(n2686), .B(n265), .Z(n2039) );
  OAI21_X4 U1862 ( .B1(n2822), .B2(n339), .A(n2720), .ZN(n2686) );
  AOI222_X2 U1863 ( .A1(n3217), .A2(n448), .B1(n315), .B2(n445), .C1(n370), 
        .C2(n442), .ZN(n2720) );
  XOR2_X2 U1864 ( .A(n2687), .B(n265), .Z(n2040) );
  OAI21_X4 U1865 ( .B1(n2823), .B2(n339), .A(n2721), .ZN(n2687) );
  AOI222_X2 U1866 ( .A1(n3217), .A2(n445), .B1(n315), .B2(n442), .C1(n370), 
        .C2(n439), .ZN(n2721) );
  XOR2_X2 U1867 ( .A(n2688), .B(n265), .Z(n2041) );
  OAI21_X4 U1868 ( .B1(n2824), .B2(n339), .A(n2722), .ZN(n2688) );
  AOI222_X2 U1869 ( .A1(n3217), .A2(n442), .B1(n315), .B2(n439), .C1(n370), 
        .C2(n436), .ZN(n2722) );
  XOR2_X2 U1870 ( .A(n2689), .B(n265), .Z(n2042) );
  OAI21_X4 U1871 ( .B1(n2825), .B2(n339), .A(n2723), .ZN(n2689) );
  AOI222_X2 U1872 ( .A1(n3217), .A2(n439), .B1(n315), .B2(n436), .C1(n370), 
        .C2(n433), .ZN(n2723) );
  XOR2_X2 U1873 ( .A(n2690), .B(n265), .Z(n2043) );
  OAI21_X4 U1874 ( .B1(n2826), .B2(n339), .A(n2724), .ZN(n2690) );
  AOI222_X2 U1875 ( .A1(n3217), .A2(n436), .B1(n315), .B2(n433), .C1(n370), 
        .C2(n430), .ZN(n2724) );
  XOR2_X2 U1876 ( .A(n2691), .B(n265), .Z(n2044) );
  OAI21_X4 U1877 ( .B1(n2827), .B2(n339), .A(n2725), .ZN(n2691) );
  AOI222_X2 U1878 ( .A1(n3217), .A2(n433), .B1(n315), .B2(n430), .C1(n370), 
        .C2(n427), .ZN(n2725) );
  XOR2_X2 U1879 ( .A(n2692), .B(n265), .Z(n2045) );
  OAI21_X4 U1880 ( .B1(n2828), .B2(n339), .A(n2726), .ZN(n2692) );
  AOI222_X2 U1881 ( .A1(n3217), .A2(n430), .B1(n315), .B2(n427), .C1(n370), 
        .C2(n424), .ZN(n2726) );
  XOR2_X2 U1882 ( .A(n2693), .B(n265), .Z(n2046) );
  OAI21_X4 U1883 ( .B1(n2829), .B2(n339), .A(n2727), .ZN(n2693) );
  AOI222_X2 U1884 ( .A1(n3217), .A2(n427), .B1(n315), .B2(n424), .C1(n370), 
        .C2(n421), .ZN(n2727) );
  XOR2_X2 U1885 ( .A(n2694), .B(n265), .Z(n2047) );
  OAI21_X4 U1886 ( .B1(n2830), .B2(n339), .A(n2728), .ZN(n2694) );
  AOI222_X2 U1887 ( .A1(n3217), .A2(n424), .B1(n315), .B2(n421), .C1(n370), 
        .C2(n418), .ZN(n2728) );
  XOR2_X2 U1888 ( .A(n2695), .B(n265), .Z(n2048) );
  OAI21_X4 U1889 ( .B1(n2831), .B2(n339), .A(n2729), .ZN(n2695) );
  AOI222_X2 U1890 ( .A1(n3217), .A2(n421), .B1(n315), .B2(n418), .C1(n370), 
        .C2(n415), .ZN(n2729) );
  XOR2_X2 U1891 ( .A(n2696), .B(n265), .Z(n2049) );
  OAI21_X4 U1892 ( .B1(n2832), .B2(n339), .A(n2730), .ZN(n2696) );
  AOI222_X2 U1893 ( .A1(n3217), .A2(n418), .B1(n315), .B2(n415), .C1(n370), 
        .C2(n412), .ZN(n2730) );
  XOR2_X2 U1894 ( .A(n2697), .B(n265), .Z(n2050) );
  OAI21_X4 U1895 ( .B1(n2833), .B2(n339), .A(n2731), .ZN(n2697) );
  AOI222_X2 U1896 ( .A1(n3217), .A2(n415), .B1(n315), .B2(n412), .C1(n370), 
        .C2(n409), .ZN(n2731) );
  XOR2_X2 U1897 ( .A(n2698), .B(n265), .Z(n2051) );
  OAI21_X4 U1898 ( .B1(n2834), .B2(n339), .A(n2732), .ZN(n2698) );
  AOI222_X2 U1899 ( .A1(n3217), .A2(n412), .B1(n315), .B2(n409), .C1(n370), 
        .C2(n406), .ZN(n2732) );
  XOR2_X2 U1900 ( .A(n2699), .B(n265), .Z(n2052) );
  OAI21_X4 U1901 ( .B1(n2835), .B2(n339), .A(n2733), .ZN(n2699) );
  AOI222_X2 U1902 ( .A1(n3217), .A2(n409), .B1(n315), .B2(n406), .C1(n370), 
        .C2(n403), .ZN(n2733) );
  XOR2_X2 U1903 ( .A(n2700), .B(n265), .Z(n2053) );
  OAI21_X4 U1904 ( .B1(n2836), .B2(n339), .A(n2734), .ZN(n2700) );
  AOI222_X2 U1905 ( .A1(n3217), .A2(n406), .B1(n315), .B2(n403), .C1(n370), 
        .C2(n400), .ZN(n2734) );
  XOR2_X2 U1906 ( .A(n2701), .B(n265), .Z(n2054) );
  OAI21_X4 U1907 ( .B1(n2837), .B2(n339), .A(n2735), .ZN(n2701) );
  AOI222_X2 U1908 ( .A1(n3217), .A2(n403), .B1(n315), .B2(n400), .C1(n370), 
        .C2(n397), .ZN(n2735) );
  XOR2_X2 U1909 ( .A(n2702), .B(n265), .Z(n2055) );
  OAI21_X4 U1910 ( .B1(n2838), .B2(n339), .A(n2736), .ZN(n2702) );
  AOI222_X2 U1911 ( .A1(n3217), .A2(n400), .B1(n315), .B2(n397), .C1(n370), 
        .C2(n393), .ZN(n2736) );
  XOR2_X2 U1912 ( .A(n2703), .B(n265), .Z(n2056) );
  OAI21_X4 U1913 ( .B1(n2839), .B2(n339), .A(n2737), .ZN(n2703) );
  AOI222_X2 U1914 ( .A1(n3217), .A2(n397), .B1(n315), .B2(n393), .C1(n370), 
        .C2(n390), .ZN(n2737) );
  XOR2_X2 U1915 ( .A(n2704), .B(n265), .Z(n2057) );
  OAI21_X4 U1916 ( .B1(n2840), .B2(n339), .A(n2738), .ZN(n2704) );
  XOR2_X2 U1918 ( .A(n2705), .B(n265), .Z(n2058) );
  AND2_X4 U1921 ( .A1(n3217), .A2(n390), .ZN(n1403) );
  XOR2_X2 U1923 ( .A(n2740), .B(n262), .Z(n2060) );
  OAI21_X4 U1924 ( .B1(n2808), .B2(n336), .A(n2774), .ZN(n2740) );
  NAND2_X4 U1925 ( .A1(n368), .A2(n484), .ZN(n2774) );
  XOR2_X2 U1926 ( .A(n2741), .B(n262), .Z(n2061) );
  OAI21_X4 U1927 ( .B1(n2809), .B2(n336), .A(n2775), .ZN(n2741) );
  AOI21_X4 U1928 ( .B1(n368), .B2(n481), .A(n1404), .ZN(n2775) );
  AND2_X4 U1929 ( .A1(n313), .A2(n484), .ZN(n1404) );
  XOR2_X2 U1930 ( .A(n2742), .B(n262), .Z(n2062) );
  OAI21_X4 U1931 ( .B1(n2810), .B2(n336), .A(n2776), .ZN(n2742) );
  AOI222_X2 U1932 ( .A1(n3152), .A2(n484), .B1(n313), .B2(n481), .C1(n368), 
        .C2(n478), .ZN(n2776) );
  XOR2_X2 U1933 ( .A(n2743), .B(n262), .Z(n2063) );
  OAI21_X4 U1934 ( .B1(n2811), .B2(n336), .A(n2777), .ZN(n2743) );
  AOI222_X2 U1935 ( .A1(n3152), .A2(n481), .B1(n313), .B2(n478), .C1(n368), 
        .C2(n475), .ZN(n2777) );
  XOR2_X2 U1936 ( .A(n2744), .B(n262), .Z(n2064) );
  OAI21_X4 U1937 ( .B1(n2812), .B2(n336), .A(n2778), .ZN(n2744) );
  AOI222_X2 U1938 ( .A1(n3151), .A2(n478), .B1(n313), .B2(n475), .C1(n368), 
        .C2(n472), .ZN(n2778) );
  XOR2_X2 U1939 ( .A(n2745), .B(n262), .Z(n2065) );
  OAI21_X4 U1940 ( .B1(n2813), .B2(n336), .A(n2779), .ZN(n2745) );
  AOI222_X2 U1941 ( .A1(n3151), .A2(n475), .B1(n313), .B2(n472), .C1(n368), 
        .C2(n469), .ZN(n2779) );
  XOR2_X2 U1942 ( .A(n2746), .B(n262), .Z(n2066) );
  OAI21_X4 U1943 ( .B1(n2814), .B2(n336), .A(n2780), .ZN(n2746) );
  AOI222_X2 U1944 ( .A1(n3151), .A2(n472), .B1(n313), .B2(n469), .C1(n368), 
        .C2(n466), .ZN(n2780) );
  XOR2_X2 U1945 ( .A(n2747), .B(n262), .Z(n2067) );
  OAI21_X4 U1946 ( .B1(n2815), .B2(n336), .A(n2781), .ZN(n2747) );
  AOI222_X2 U1947 ( .A1(n3152), .A2(n469), .B1(n313), .B2(n466), .C1(n368), 
        .C2(n463), .ZN(n2781) );
  XOR2_X2 U1948 ( .A(n2748), .B(n262), .Z(n2068) );
  OAI21_X4 U1949 ( .B1(n2816), .B2(n336), .A(n2782), .ZN(n2748) );
  AOI222_X2 U1950 ( .A1(n3152), .A2(n466), .B1(n313), .B2(n463), .C1(n368), 
        .C2(n460), .ZN(n2782) );
  XOR2_X2 U1951 ( .A(n2749), .B(n262), .Z(n2069) );
  OAI21_X4 U1952 ( .B1(n2817), .B2(n336), .A(n2783), .ZN(n2749) );
  AOI222_X2 U1953 ( .A1(n3151), .A2(n463), .B1(n313), .B2(n460), .C1(n368), 
        .C2(n457), .ZN(n2783) );
  XOR2_X2 U1954 ( .A(n2750), .B(n262), .Z(n2070) );
  OAI21_X4 U1955 ( .B1(n2818), .B2(n336), .A(n2784), .ZN(n2750) );
  AOI222_X2 U1956 ( .A1(n3152), .A2(n460), .B1(n313), .B2(n457), .C1(n368), 
        .C2(n454), .ZN(n2784) );
  XOR2_X2 U1957 ( .A(n2751), .B(n262), .Z(n2071) );
  OAI21_X4 U1958 ( .B1(n2819), .B2(n336), .A(n2785), .ZN(n2751) );
  AOI222_X2 U1959 ( .A1(n3151), .A2(n457), .B1(n313), .B2(n454), .C1(n368), 
        .C2(n451), .ZN(n2785) );
  XOR2_X2 U1960 ( .A(n2752), .B(n262), .Z(n2072) );
  OAI21_X4 U1961 ( .B1(n2820), .B2(n336), .A(n2786), .ZN(n2752) );
  AOI222_X2 U1962 ( .A1(n3152), .A2(n454), .B1(n313), .B2(n451), .C1(n368), 
        .C2(n448), .ZN(n2786) );
  XOR2_X2 U1963 ( .A(n2753), .B(n262), .Z(n2073) );
  OAI21_X4 U1964 ( .B1(n2821), .B2(n336), .A(n2787), .ZN(n2753) );
  AOI222_X2 U1965 ( .A1(n3151), .A2(n451), .B1(n313), .B2(n448), .C1(n368), 
        .C2(n445), .ZN(n2787) );
  XOR2_X2 U1966 ( .A(n2754), .B(n262), .Z(n2074) );
  OAI21_X4 U1967 ( .B1(n2822), .B2(n336), .A(n2788), .ZN(n2754) );
  AOI222_X2 U1968 ( .A1(n3152), .A2(n448), .B1(n313), .B2(n445), .C1(n368), 
        .C2(n442), .ZN(n2788) );
  XOR2_X2 U1969 ( .A(n2755), .B(n262), .Z(n2075) );
  OAI21_X4 U1970 ( .B1(n2823), .B2(n336), .A(n2789), .ZN(n2755) );
  AOI222_X2 U1971 ( .A1(n3151), .A2(n445), .B1(n313), .B2(n442), .C1(n368), 
        .C2(n439), .ZN(n2789) );
  XOR2_X2 U1972 ( .A(n2756), .B(n262), .Z(n2076) );
  OAI21_X4 U1973 ( .B1(n2824), .B2(n336), .A(n2790), .ZN(n2756) );
  AOI222_X2 U1974 ( .A1(n3152), .A2(n442), .B1(n313), .B2(n439), .C1(n368), 
        .C2(n436), .ZN(n2790) );
  XOR2_X2 U1975 ( .A(n2757), .B(n262), .Z(n2077) );
  OAI21_X4 U1976 ( .B1(n2825), .B2(n336), .A(n2791), .ZN(n2757) );
  AOI222_X2 U1977 ( .A1(n3152), .A2(n439), .B1(n313), .B2(n436), .C1(n368), 
        .C2(n433), .ZN(n2791) );
  XOR2_X2 U1978 ( .A(n2758), .B(n262), .Z(n2078) );
  OAI21_X4 U1979 ( .B1(n2826), .B2(n336), .A(n2792), .ZN(n2758) );
  AOI222_X2 U1980 ( .A1(n3151), .A2(n436), .B1(n313), .B2(n433), .C1(n368), 
        .C2(n430), .ZN(n2792) );
  XOR2_X2 U1981 ( .A(n2759), .B(n262), .Z(n2079) );
  OAI21_X4 U1982 ( .B1(n2827), .B2(n336), .A(n2793), .ZN(n2759) );
  AOI222_X2 U1983 ( .A1(n3152), .A2(n433), .B1(n313), .B2(n430), .C1(n368), 
        .C2(n427), .ZN(n2793) );
  XOR2_X2 U1984 ( .A(n2760), .B(n262), .Z(n2080) );
  OAI21_X4 U1985 ( .B1(n2828), .B2(n336), .A(n2794), .ZN(n2760) );
  AOI222_X2 U1986 ( .A1(n3151), .A2(n430), .B1(n313), .B2(n427), .C1(n368), 
        .C2(n424), .ZN(n2794) );
  XOR2_X2 U1987 ( .A(n2761), .B(n262), .Z(n2081) );
  OAI21_X4 U1988 ( .B1(n2829), .B2(n336), .A(n2795), .ZN(n2761) );
  AOI222_X2 U1989 ( .A1(n3151), .A2(n427), .B1(n313), .B2(n424), .C1(n368), 
        .C2(n421), .ZN(n2795) );
  XOR2_X2 U1990 ( .A(n2762), .B(n262), .Z(n2082) );
  OAI21_X4 U1991 ( .B1(n2830), .B2(n336), .A(n2796), .ZN(n2762) );
  AOI222_X2 U1992 ( .A1(n3151), .A2(n424), .B1(n313), .B2(n421), .C1(n368), 
        .C2(n418), .ZN(n2796) );
  XOR2_X2 U1993 ( .A(n2763), .B(n262), .Z(n2083) );
  OAI21_X4 U1994 ( .B1(n2831), .B2(n336), .A(n2797), .ZN(n2763) );
  AOI222_X2 U1995 ( .A1(n3151), .A2(n421), .B1(n313), .B2(n418), .C1(n368), 
        .C2(n415), .ZN(n2797) );
  XOR2_X2 U1996 ( .A(n2764), .B(n262), .Z(n2084) );
  OAI21_X4 U1997 ( .B1(n2832), .B2(n336), .A(n2798), .ZN(n2764) );
  AOI222_X2 U1998 ( .A1(n3152), .A2(n418), .B1(n313), .B2(n415), .C1(n368), 
        .C2(n412), .ZN(n2798) );
  XOR2_X2 U1999 ( .A(n2765), .B(n262), .Z(n2085) );
  OAI21_X4 U2000 ( .B1(n2833), .B2(n336), .A(n2799), .ZN(n2765) );
  AOI222_X2 U2001 ( .A1(n3152), .A2(n415), .B1(n313), .B2(n412), .C1(n368), 
        .C2(n409), .ZN(n2799) );
  XOR2_X2 U2002 ( .A(n2766), .B(n262), .Z(n2086) );
  OAI21_X4 U2003 ( .B1(n2834), .B2(n336), .A(n2800), .ZN(n2766) );
  AOI222_X2 U2004 ( .A1(n3151), .A2(n412), .B1(n313), .B2(n409), .C1(n368), 
        .C2(n406), .ZN(n2800) );
  XOR2_X2 U2005 ( .A(n2767), .B(n262), .Z(n2087) );
  OAI21_X4 U2006 ( .B1(n2835), .B2(n336), .A(n2801), .ZN(n2767) );
  AOI222_X2 U2007 ( .A1(n3152), .A2(n409), .B1(n313), .B2(n406), .C1(n368), 
        .C2(n403), .ZN(n2801) );
  XOR2_X2 U2008 ( .A(n2768), .B(n262), .Z(n2088) );
  OAI21_X4 U2009 ( .B1(n2836), .B2(n336), .A(n2802), .ZN(n2768) );
  AOI222_X2 U2010 ( .A1(n3151), .A2(n406), .B1(n313), .B2(n403), .C1(n368), 
        .C2(n400), .ZN(n2802) );
  XOR2_X2 U2011 ( .A(n2769), .B(n262), .Z(n2089) );
  OAI21_X4 U2012 ( .B1(n2837), .B2(n336), .A(n2803), .ZN(n2769) );
  AOI222_X2 U2013 ( .A1(n3152), .A2(n403), .B1(n313), .B2(n400), .C1(n368), 
        .C2(n397), .ZN(n2803) );
  XOR2_X2 U2014 ( .A(n2770), .B(n262), .Z(n2090) );
  OAI21_X4 U2015 ( .B1(n2838), .B2(n336), .A(n2804), .ZN(n2770) );
  AOI222_X2 U2016 ( .A1(n3152), .A2(n400), .B1(n313), .B2(n397), .C1(n368), 
        .C2(n393), .ZN(n2804) );
  XOR2_X2 U2017 ( .A(n2771), .B(n262), .Z(n2091) );
  OAI21_X4 U2018 ( .B1(n2839), .B2(n336), .A(n2805), .ZN(n2771) );
  AOI222_X2 U2019 ( .A1(n3151), .A2(n397), .B1(n313), .B2(n393), .C1(n368), 
        .C2(n390), .ZN(n2805) );
  XOR2_X2 U2020 ( .A(n2772), .B(n262), .Z(n678) );
  OAI21_X4 U2021 ( .B1(n2840), .B2(n336), .A(n2806), .ZN(n2772) );
  AND2_X4 U2026 ( .A1(n3151), .A2(n390), .ZN(n1406) );
  AND3_X4 U2103 ( .A1(n2908), .A2(n2919), .A3(a[31]), .ZN(n388) );
  AND3_X4 U2107 ( .A1(n2931), .A2(n2909), .A3(n2920), .ZN(n386) );
  AND3_X4 U2112 ( .A1(n2932), .A2(n2910), .A3(n2921), .ZN(n384) );
  AND3_X4 U2117 ( .A1(n2933), .A2(n2911), .A3(n2922), .ZN(n382) );
  AND3_X4 U2122 ( .A1(n2934), .A2(n2912), .A3(n2923), .ZN(n380) );
  AND3_X4 U2127 ( .A1(n2935), .A2(n2913), .A3(n2924), .ZN(n378) );
  AND3_X4 U2132 ( .A1(n2936), .A2(n2914), .A3(n2925), .ZN(n376) );
  AND3_X4 U2137 ( .A1(n2937), .A2(n2915), .A3(n2926), .ZN(n374) );
  XNOR2_X2 U2140 ( .A(n268), .B(a[9]), .ZN(n2915) );
  XOR2_X2 U2141 ( .A(a[10]), .B(n271), .Z(n2937) );
  AND3_X4 U2142 ( .A1(n2938), .A2(n2916), .A3(n2927), .ZN(n372) );
  XNOR2_X2 U2145 ( .A(n265), .B(a[6]), .ZN(n2916) );
  XOR2_X2 U2146 ( .A(a[7]), .B(n268), .Z(n2938) );
  AND3_X4 U2147 ( .A1(n2939), .A2(n2917), .A3(n2928), .ZN(n370) );
  XNOR2_X2 U2150 ( .A(n262), .B(a[3]), .ZN(n2917) );
  AND3_X4 U2152 ( .A1(n2940), .A2(n2929), .A3(n2918), .ZN(n368) );
  XNOR2_X2 U2158 ( .A(n1441), .B(n1440), .ZN(n2843) );
  NAND2_X4 U2159 ( .A1(n1441), .A2(n484), .ZN(n2808) );
  XOR2_X2 U2162 ( .A(n1452), .B(n1407), .Z(n2844) );
  OAI21_X4 U2163 ( .B1(n1600), .B2(n1442), .A(n1443), .ZN(n1441) );
  NAND2_X4 U2164 ( .A1(n1528), .A2(n1444), .ZN(n1442) );
  AOI21_X4 U2165 ( .B1(n1529), .B2(n1444), .A(n1445), .ZN(n1443) );
  NOR2_X4 U2166 ( .A1(n1488), .A2(n1446), .ZN(n1444) );
  OAI21_X4 U2167 ( .B1(n1489), .B2(n1446), .A(n1447), .ZN(n1445) );
  NAND2_X4 U2168 ( .A1(n1468), .A2(n1448), .ZN(n1446) );
  AOI21_X4 U2169 ( .B1(n1448), .B2(n1469), .A(n1449), .ZN(n1447) );
  NOR2_X4 U2170 ( .A1(n1459), .A2(n1450), .ZN(n1448) );
  OAI21_X4 U2171 ( .B1(n1450), .B2(n1462), .A(n1451), .ZN(n1449) );
  NAND2_X4 U2172 ( .A1(n1689), .A2(n1451), .ZN(n1407) );
  NOR2_X4 U2174 ( .A1(n481), .A2(n484), .ZN(n1450) );
  NAND2_X4 U2175 ( .A1(n481), .A2(n484), .ZN(n1451) );
  XOR2_X2 U2176 ( .A(n1463), .B(n1408), .Z(n2845) );
  AOI21_X4 U2177 ( .B1(n1599), .B2(n1453), .A(n1454), .ZN(n1452) );
  NOR2_X4 U2178 ( .A1(n1530), .A2(n1455), .ZN(n1453) );
  OAI21_X4 U2179 ( .B1(n1531), .B2(n1455), .A(n1456), .ZN(n1454) );
  NAND2_X4 U2180 ( .A1(n1457), .A2(n1490), .ZN(n1455) );
  AOI21_X4 U2181 ( .B1(n1457), .B2(n1491), .A(n1458), .ZN(n1456) );
  NOR2_X4 U2182 ( .A1(n1470), .A2(n1459), .ZN(n1457) );
  OAI21_X4 U2183 ( .B1(n1471), .B2(n1459), .A(n1462), .ZN(n1458) );
  NAND2_X4 U2186 ( .A1(n1690), .A2(n1462), .ZN(n1408) );
  NOR2_X4 U2188 ( .A1(n478), .A2(n481), .ZN(n1459) );
  NAND2_X4 U2189 ( .A1(n478), .A2(n481), .ZN(n1462) );
  XOR2_X2 U2190 ( .A(n1476), .B(n1409), .Z(n2846) );
  AOI21_X4 U2191 ( .B1(n1599), .B2(n1464), .A(n1465), .ZN(n1463) );
  NOR2_X4 U2192 ( .A1(n1530), .A2(n1466), .ZN(n1464) );
  OAI21_X4 U2193 ( .B1(n1531), .B2(n1466), .A(n1467), .ZN(n1465) );
  NAND2_X4 U2194 ( .A1(n1490), .A2(n1468), .ZN(n1466) );
  AOI21_X4 U2195 ( .B1(n1491), .B2(n1468), .A(n1469), .ZN(n1467) );
  NOR2_X4 U2200 ( .A1(n1483), .A2(n1474), .ZN(n1468) );
  OAI21_X4 U2201 ( .B1(n1474), .B2(n1484), .A(n1475), .ZN(n1469) );
  NAND2_X4 U2202 ( .A1(n1691), .A2(n1475), .ZN(n1409) );
  NOR2_X4 U2204 ( .A1(n475), .A2(n478), .ZN(n1474) );
  NAND2_X4 U2205 ( .A1(n475), .A2(n478), .ZN(n1475) );
  XOR2_X2 U2206 ( .A(n1485), .B(n1410), .Z(n2847) );
  AOI21_X4 U2207 ( .B1(n1599), .B2(n1477), .A(n1478), .ZN(n1476) );
  NOR2_X4 U2208 ( .A1(n1530), .A2(n1479), .ZN(n1477) );
  OAI21_X4 U2209 ( .B1(n1531), .B2(n1479), .A(n1480), .ZN(n1478) );
  NAND2_X4 U2210 ( .A1(n1490), .A2(n1692), .ZN(n1479) );
  AOI21_X4 U2211 ( .B1(n1491), .B2(n1692), .A(n1482), .ZN(n1480) );
  NAND2_X4 U2214 ( .A1(n1692), .A2(n1484), .ZN(n1410) );
  NOR2_X4 U2216 ( .A1(n472), .A2(n475), .ZN(n1483) );
  NAND2_X4 U2217 ( .A1(n472), .A2(n475), .ZN(n1484) );
  XOR2_X2 U2218 ( .A(n1498), .B(n1411), .Z(n2848) );
  AOI21_X4 U2219 ( .B1(n1599), .B2(n1486), .A(n1487), .ZN(n1485) );
  NOR2_X4 U2220 ( .A1(n1530), .A2(n1488), .ZN(n1486) );
  OAI21_X4 U2221 ( .B1(n1531), .B2(n1488), .A(n1489), .ZN(n1487) );
  NAND2_X4 U2226 ( .A1(n1512), .A2(n1494), .ZN(n1488) );
  AOI21_X4 U2227 ( .B1(n1494), .B2(n1513), .A(n1495), .ZN(n1489) );
  NOR2_X4 U2228 ( .A1(n1505), .A2(n1496), .ZN(n1494) );
  OAI21_X4 U2229 ( .B1(n1496), .B2(n1506), .A(n1497), .ZN(n1495) );
  NAND2_X4 U2230 ( .A1(n1693), .A2(n1497), .ZN(n1411) );
  NOR2_X4 U2232 ( .A1(n469), .A2(n472), .ZN(n1496) );
  NAND2_X4 U2233 ( .A1(n469), .A2(n472), .ZN(n1497) );
  XOR2_X2 U2234 ( .A(n1507), .B(n1412), .Z(n2849) );
  AOI21_X4 U2235 ( .B1(n1599), .B2(n1499), .A(n1500), .ZN(n1498) );
  NOR2_X4 U2236 ( .A1(n1530), .A2(n1501), .ZN(n1499) );
  OAI21_X4 U2237 ( .B1(n1531), .B2(n1501), .A(n1502), .ZN(n1500) );
  NAND2_X4 U2238 ( .A1(n1512), .A2(n1694), .ZN(n1501) );
  AOI21_X4 U2239 ( .B1(n1513), .B2(n1694), .A(n1504), .ZN(n1502) );
  NAND2_X4 U2242 ( .A1(n1694), .A2(n1506), .ZN(n1412) );
  NOR2_X4 U2244 ( .A1(n466), .A2(n469), .ZN(n1505) );
  NAND2_X4 U2245 ( .A1(n466), .A2(n469), .ZN(n1506) );
  XOR2_X2 U2246 ( .A(n1520), .B(n1413), .Z(n2850) );
  AOI21_X4 U2247 ( .B1(n1599), .B2(n1508), .A(n1509), .ZN(n1507) );
  NOR2_X4 U2248 ( .A1(n1530), .A2(n1510), .ZN(n1508) );
  OAI21_X4 U2249 ( .B1(n1531), .B2(n1510), .A(n1511), .ZN(n1509) );
  NOR2_X4 U2256 ( .A1(n1523), .A2(n1518), .ZN(n1512) );
  OAI21_X4 U2257 ( .B1(n1518), .B2(n1526), .A(n1519), .ZN(n1513) );
  NAND2_X4 U2258 ( .A1(n1695), .A2(n1519), .ZN(n1413) );
  NOR2_X4 U2260 ( .A1(n463), .A2(n466), .ZN(n1518) );
  NAND2_X4 U2261 ( .A1(n463), .A2(n466), .ZN(n1519) );
  XOR2_X2 U2262 ( .A(n1527), .B(n1414), .Z(n2851) );
  AOI21_X4 U2263 ( .B1(n1599), .B2(n1521), .A(n1522), .ZN(n1520) );
  NOR2_X4 U2264 ( .A1(n1530), .A2(n1523), .ZN(n1521) );
  OAI21_X4 U2265 ( .B1(n1531), .B2(n1523), .A(n1526), .ZN(n1522) );
  NAND2_X4 U2268 ( .A1(n1696), .A2(n1526), .ZN(n1414) );
  NOR2_X4 U2270 ( .A1(n460), .A2(n463), .ZN(n1523) );
  NAND2_X4 U2271 ( .A1(n460), .A2(n463), .ZN(n1526) );
  XOR2_X2 U2272 ( .A(n1540), .B(n1415), .Z(n2852) );
  AOI21_X4 U2273 ( .B1(n1599), .B2(n1528), .A(n1529), .ZN(n1527) );
  NOR2_X4 U2278 ( .A1(n1568), .A2(n1534), .ZN(n1528) );
  OAI21_X4 U2279 ( .B1(n1569), .B2(n1534), .A(n1535), .ZN(n1529) );
  NAND2_X4 U2280 ( .A1(n1552), .A2(n1536), .ZN(n1534) );
  AOI21_X4 U2281 ( .B1(n1536), .B2(n1555), .A(n1537), .ZN(n1535) );
  NOR2_X4 U2282 ( .A1(n1543), .A2(n1538), .ZN(n1536) );
  OAI21_X4 U2283 ( .B1(n1538), .B2(n1546), .A(n1539), .ZN(n1537) );
  NAND2_X4 U2284 ( .A1(n1697), .A2(n1539), .ZN(n1415) );
  NOR2_X4 U2286 ( .A1(n457), .A2(n460), .ZN(n1538) );
  NAND2_X4 U2287 ( .A1(n457), .A2(n460), .ZN(n1539) );
  XOR2_X2 U2288 ( .A(n1547), .B(n1416), .Z(n2853) );
  AOI21_X4 U2289 ( .B1(n1599), .B2(n1541), .A(n1542), .ZN(n1540) );
  NOR2_X4 U2290 ( .A1(n1550), .A2(n1543), .ZN(n1541) );
  OAI21_X4 U2291 ( .B1(n1551), .B2(n1543), .A(n1546), .ZN(n1542) );
  NAND2_X4 U2294 ( .A1(n1698), .A2(n1546), .ZN(n1416) );
  NOR2_X4 U2296 ( .A1(n454), .A2(n457), .ZN(n1543) );
  NAND2_X4 U2297 ( .A1(n454), .A2(n457), .ZN(n1546) );
  XOR2_X2 U2298 ( .A(n1558), .B(n1417), .Z(n2854) );
  AOI21_X4 U2299 ( .B1(n1599), .B2(n1548), .A(n1549), .ZN(n1547) );
  NAND2_X4 U2302 ( .A1(n1570), .A2(n1552), .ZN(n1550) );
  AOI21_X4 U2303 ( .B1(n1571), .B2(n1552), .A(n1555), .ZN(n1551) );
  NOR2_X4 U2306 ( .A1(n1561), .A2(n1556), .ZN(n1552) );
  OAI21_X4 U2307 ( .B1(n1556), .B2(n1564), .A(n1557), .ZN(n1555) );
  NAND2_X4 U2308 ( .A1(n1699), .A2(n1557), .ZN(n1417) );
  NOR2_X4 U2310 ( .A1(n451), .A2(n454), .ZN(n1556) );
  NAND2_X4 U2311 ( .A1(n451), .A2(n454), .ZN(n1557) );
  XOR2_X2 U2312 ( .A(n1565), .B(n1418), .Z(n2855) );
  AOI21_X4 U2313 ( .B1(n1599), .B2(n1559), .A(n1560), .ZN(n1558) );
  NOR2_X4 U2314 ( .A1(n1568), .A2(n1561), .ZN(n1559) );
  OAI21_X4 U2315 ( .B1(n1569), .B2(n1561), .A(n1564), .ZN(n1560) );
  NAND2_X4 U2318 ( .A1(n1700), .A2(n1564), .ZN(n1418) );
  NOR2_X4 U2320 ( .A1(n448), .A2(n451), .ZN(n1561) );
  NAND2_X4 U2321 ( .A1(n448), .A2(n451), .ZN(n1564) );
  XOR2_X2 U2322 ( .A(n1578), .B(n1419), .Z(n2856) );
  AOI21_X4 U2323 ( .B1(n1599), .B2(n1570), .A(n1571), .ZN(n1565) );
  NAND2_X4 U2330 ( .A1(n1586), .A2(n1574), .ZN(n1568) );
  AOI21_X4 U2331 ( .B1(n1574), .B2(n1587), .A(n1575), .ZN(n1569) );
  NOR2_X4 U2332 ( .A1(n1581), .A2(n1576), .ZN(n1574) );
  OAI21_X4 U2333 ( .B1(n1576), .B2(n1584), .A(n1577), .ZN(n1575) );
  NAND2_X4 U2334 ( .A1(n1701), .A2(n1577), .ZN(n1419) );
  NOR2_X4 U2336 ( .A1(n445), .A2(n448), .ZN(n1576) );
  NAND2_X4 U2337 ( .A1(n445), .A2(n448), .ZN(n1577) );
  XOR2_X2 U2338 ( .A(n1585), .B(n1420), .Z(n2857) );
  AOI21_X4 U2339 ( .B1(n1599), .B2(n1579), .A(n1580), .ZN(n1578) );
  NOR2_X4 U2340 ( .A1(n1588), .A2(n1581), .ZN(n1579) );
  OAI21_X4 U2341 ( .B1(n1589), .B2(n1581), .A(n1584), .ZN(n1580) );
  NAND2_X4 U2344 ( .A1(n1702), .A2(n1584), .ZN(n1420) );
  NOR2_X4 U2346 ( .A1(n442), .A2(n445), .ZN(n1581) );
  NAND2_X4 U2347 ( .A1(n442), .A2(n445), .ZN(n1584) );
  XOR2_X2 U2348 ( .A(n1594), .B(n1421), .Z(n2858) );
  AOI21_X4 U2349 ( .B1(n1599), .B2(n1586), .A(n1587), .ZN(n1585) );
  NOR2_X4 U2354 ( .A1(n1597), .A2(n1592), .ZN(n1586) );
  OAI21_X4 U2355 ( .B1(n1592), .B2(n1598), .A(n1593), .ZN(n1587) );
  NAND2_X4 U2356 ( .A1(n1703), .A2(n1593), .ZN(n1421) );
  NOR2_X4 U2358 ( .A1(n439), .A2(n442), .ZN(n1592) );
  NAND2_X4 U2359 ( .A1(n439), .A2(n442), .ZN(n1593) );
  XNOR2_X2 U2360 ( .A(n1599), .B(n1422), .ZN(n2859) );
  AOI21_X4 U2361 ( .B1(n1599), .B2(n1704), .A(n1596), .ZN(n1594) );
  NAND2_X4 U2364 ( .A1(n1704), .A2(n1598), .ZN(n1422) );
  NOR2_X4 U2366 ( .A1(n436), .A2(n439), .ZN(n1597) );
  NAND2_X4 U2367 ( .A1(n436), .A2(n439), .ZN(n1598) );
  XOR2_X2 U2368 ( .A(n1609), .B(n1423), .Z(n2860) );
  AOI21_X4 U2370 ( .B1(n1655), .B2(n1601), .A(n1602), .ZN(n1600) );
  NOR2_X4 U2371 ( .A1(n1629), .A2(n1603), .ZN(n1601) );
  OAI21_X4 U2372 ( .B1(n1630), .B2(n1603), .A(n1604), .ZN(n1602) );
  NAND2_X4 U2373 ( .A1(n1617), .A2(n1605), .ZN(n1603) );
  AOI21_X4 U2374 ( .B1(n1605), .B2(n1620), .A(n1606), .ZN(n1604) );
  NOR2_X4 U2375 ( .A1(n1612), .A2(n1607), .ZN(n1605) );
  OAI21_X4 U2376 ( .B1(n1607), .B2(n1613), .A(n1608), .ZN(n1606) );
  NAND2_X4 U2377 ( .A1(n1705), .A2(n1608), .ZN(n1423) );
  NOR2_X4 U2379 ( .A1(n433), .A2(n436), .ZN(n1607) );
  NAND2_X4 U2380 ( .A1(n433), .A2(n436), .ZN(n1608) );
  XNOR2_X2 U2381 ( .A(n1614), .B(n1424), .ZN(n2861) );
  AOI21_X4 U2382 ( .B1(n1614), .B2(n1706), .A(n1611), .ZN(n1609) );
  NAND2_X4 U2385 ( .A1(n1706), .A2(n1613), .ZN(n1424) );
  NOR2_X4 U2387 ( .A1(n430), .A2(n433), .ZN(n1612) );
  NAND2_X4 U2388 ( .A1(n430), .A2(n433), .ZN(n1613) );
  XOR2_X2 U2389 ( .A(n1623), .B(n1425), .Z(n2862) );
  OAI21_X4 U2390 ( .B1(n1654), .B2(n1615), .A(n1616), .ZN(n1614) );
  NAND2_X4 U2391 ( .A1(n1631), .A2(n1617), .ZN(n1615) );
  AOI21_X4 U2392 ( .B1(n1632), .B2(n1617), .A(n1620), .ZN(n1616) );
  NOR2_X4 U2395 ( .A1(n1626), .A2(n1621), .ZN(n1617) );
  OAI21_X4 U2396 ( .B1(n1621), .B2(n1627), .A(n1622), .ZN(n1620) );
  NAND2_X4 U2397 ( .A1(n1707), .A2(n1622), .ZN(n1425) );
  NOR2_X4 U2399 ( .A1(n427), .A2(n430), .ZN(n1621) );
  NAND2_X4 U2400 ( .A1(n427), .A2(n430), .ZN(n1622) );
  XNOR2_X2 U2401 ( .A(n1628), .B(n1426), .ZN(n2863) );
  AOI21_X4 U2402 ( .B1(n1628), .B2(n1708), .A(n1625), .ZN(n1623) );
  NAND2_X4 U2405 ( .A1(n1708), .A2(n1627), .ZN(n1426) );
  NOR2_X4 U2407 ( .A1(n424), .A2(n427), .ZN(n1626) );
  NAND2_X4 U2408 ( .A1(n424), .A2(n427), .ZN(n1627) );
  XOR2_X2 U2409 ( .A(n1639), .B(n1427), .Z(n2864) );
  OAI21_X4 U2410 ( .B1(n1654), .B2(n1629), .A(n1630), .ZN(n1628) );
  NAND2_X4 U2415 ( .A1(n1647), .A2(n1635), .ZN(n1629) );
  AOI21_X4 U2416 ( .B1(n1635), .B2(n1648), .A(n1636), .ZN(n1630) );
  NOR2_X4 U2417 ( .A1(n1642), .A2(n1637), .ZN(n1635) );
  OAI21_X4 U2418 ( .B1(n1637), .B2(n1643), .A(n1638), .ZN(n1636) );
  NAND2_X4 U2419 ( .A1(n1709), .A2(n1638), .ZN(n1427) );
  NOR2_X4 U2421 ( .A1(n421), .A2(n424), .ZN(n1637) );
  NAND2_X4 U2422 ( .A1(n421), .A2(n424), .ZN(n1638) );
  XNOR2_X2 U2423 ( .A(n1644), .B(n1428), .ZN(n2865) );
  AOI21_X4 U2424 ( .B1(n1644), .B2(n1710), .A(n1641), .ZN(n1639) );
  NAND2_X4 U2427 ( .A1(n1710), .A2(n1643), .ZN(n1428) );
  NOR2_X4 U2429 ( .A1(n418), .A2(n421), .ZN(n1642) );
  NAND2_X4 U2430 ( .A1(n418), .A2(n421), .ZN(n1643) );
  XNOR2_X2 U2431 ( .A(n1651), .B(n1429), .ZN(n2866) );
  OAI21_X4 U2432 ( .B1(n1654), .B2(n1645), .A(n1646), .ZN(n1644) );
  NOR2_X4 U2435 ( .A1(n1652), .A2(n1649), .ZN(n1647) );
  OAI21_X4 U2436 ( .B1(n1649), .B2(n1653), .A(n1650), .ZN(n1648) );
  NAND2_X4 U2437 ( .A1(n1711), .A2(n1650), .ZN(n1429) );
  NOR2_X4 U2439 ( .A1(n415), .A2(n418), .ZN(n1649) );
  NAND2_X4 U2440 ( .A1(n415), .A2(n418), .ZN(n1650) );
  XOR2_X2 U2441 ( .A(n1654), .B(n1430), .Z(n2867) );
  OAI21_X4 U2442 ( .B1(n1654), .B2(n1652), .A(n1653), .ZN(n1651) );
  NAND2_X4 U2443 ( .A1(n1712), .A2(n1653), .ZN(n1430) );
  NOR2_X4 U2445 ( .A1(n412), .A2(n415), .ZN(n1652) );
  NAND2_X4 U2446 ( .A1(n412), .A2(n415), .ZN(n1653) );
  XNOR2_X2 U2447 ( .A(n1662), .B(n1431), .ZN(n2868) );
  OAI21_X4 U2449 ( .B1(n1676), .B2(n1656), .A(n1657), .ZN(n1655) );
  NAND2_X4 U2450 ( .A1(n1666), .A2(n1658), .ZN(n1656) );
  AOI21_X4 U2451 ( .B1(n1658), .B2(n1667), .A(n1659), .ZN(n1657) );
  NOR2_X4 U2452 ( .A1(n1663), .A2(n1660), .ZN(n1658) );
  OAI21_X4 U2453 ( .B1(n1660), .B2(n1664), .A(n1661), .ZN(n1659) );
  NAND2_X4 U2454 ( .A1(n1713), .A2(n1661), .ZN(n1431) );
  NOR2_X4 U2456 ( .A1(n409), .A2(n412), .ZN(n1660) );
  NAND2_X4 U2457 ( .A1(n409), .A2(n412), .ZN(n1661) );
  XOR2_X2 U2458 ( .A(n1665), .B(n1432), .Z(n2869) );
  OAI21_X4 U2459 ( .B1(n1665), .B2(n1663), .A(n1664), .ZN(n1662) );
  NAND2_X4 U2460 ( .A1(n1714), .A2(n1664), .ZN(n1432) );
  NOR2_X4 U2462 ( .A1(n406), .A2(n409), .ZN(n1663) );
  NAND2_X4 U2463 ( .A1(n406), .A2(n409), .ZN(n1664) );
  XOR2_X2 U2464 ( .A(n1670), .B(n1433), .Z(n2870) );
  AOI21_X4 U2465 ( .B1(n1675), .B2(n1666), .A(n1667), .ZN(n1665) );
  NOR2_X4 U2466 ( .A1(n1673), .A2(n1668), .ZN(n1666) );
  OAI21_X4 U2467 ( .B1(n1668), .B2(n1674), .A(n1669), .ZN(n1667) );
  NAND2_X4 U2468 ( .A1(n1715), .A2(n1669), .ZN(n1433) );
  NOR2_X4 U2470 ( .A1(n403), .A2(n406), .ZN(n1668) );
  NAND2_X4 U2471 ( .A1(n403), .A2(n406), .ZN(n1669) );
  XNOR2_X2 U2472 ( .A(n1675), .B(n1434), .ZN(n2871) );
  AOI21_X4 U2473 ( .B1(n1675), .B2(n1716), .A(n1672), .ZN(n1670) );
  NAND2_X4 U2476 ( .A1(n1716), .A2(n1674), .ZN(n1434) );
  NOR2_X4 U2478 ( .A1(n400), .A2(n403), .ZN(n1673) );
  NAND2_X4 U2479 ( .A1(n400), .A2(n403), .ZN(n1674) );
  XNOR2_X2 U2480 ( .A(n1681), .B(n1435), .ZN(n2872) );
  AOI21_X4 U2482 ( .B1(n1677), .B2(n1685), .A(n1678), .ZN(n1676) );
  NOR2_X4 U2483 ( .A1(n1682), .A2(n1679), .ZN(n1677) );
  OAI21_X4 U2484 ( .B1(n1679), .B2(n1683), .A(n1680), .ZN(n1678) );
  NAND2_X4 U2485 ( .A1(n1717), .A2(n1680), .ZN(n1435) );
  NOR2_X4 U2487 ( .A1(n397), .A2(n400), .ZN(n1679) );
  NAND2_X4 U2488 ( .A1(n397), .A2(n400), .ZN(n1680) );
  XOR2_X2 U2489 ( .A(n1436), .B(n1684), .Z(n2873) );
  OAI21_X4 U2490 ( .B1(n1682), .B2(n1684), .A(n1683), .ZN(n1681) );
  NAND2_X4 U2491 ( .A1(n1718), .A2(n1683), .ZN(n1436) );
  NOR2_X4 U2493 ( .A1(n393), .A2(n397), .ZN(n1682) );
  NAND2_X4 U2494 ( .A1(n393), .A2(n397), .ZN(n1683) );
  NAND2_X4 U2498 ( .A1(n1719), .A2(n1684), .ZN(n2840) );
  NOR2_X4 U2500 ( .A1(n390), .A2(n393), .ZN(n1686) );
  NAND2_X4 U2501 ( .A1(n390), .A2(n393), .ZN(n1684) );
  XOR2_X1 U2506 ( .A(a[28]), .B(n289), .Z(n2931) );
  XNOR2_X1 U2507 ( .A(a[27]), .B(a[28]), .ZN(n2920) );
  XOR2_X1 U2508 ( .A(a[25]), .B(n286), .Z(n2932) );
  XNOR2_X1 U2509 ( .A(a[24]), .B(a[25]), .ZN(n2921) );
  XOR2_X1 U2510 ( .A(a[22]), .B(n283), .Z(n2933) );
  XNOR2_X1 U2511 ( .A(n280), .B(a[21]), .ZN(n2911) );
  XNOR2_X1 U2512 ( .A(a[21]), .B(a[22]), .ZN(n2922) );
  XOR2_X1 U2513 ( .A(a[19]), .B(n280), .Z(n2934) );
  XNOR2_X1 U2514 ( .A(n277), .B(a[18]), .ZN(n2912) );
  XNOR2_X1 U2515 ( .A(a[18]), .B(a[19]), .ZN(n2923) );
  XOR2_X1 U2516 ( .A(a[16]), .B(n277), .Z(n2935) );
  XNOR2_X1 U2517 ( .A(n274), .B(a[15]), .ZN(n2913) );
  XNOR2_X1 U2518 ( .A(a[15]), .B(a[16]), .ZN(n2924) );
  XOR2_X1 U2519 ( .A(a[13]), .B(n274), .Z(n2936) );
  XNOR2_X1 U2520 ( .A(n271), .B(a[12]), .ZN(n2914) );
  XNOR2_X1 U2521 ( .A(a[12]), .B(a[13]), .ZN(n2925) );
  XNOR2_X1 U2522 ( .A(a[9]), .B(a[10]), .ZN(n2926) );
  XNOR2_X1 U2523 ( .A(a[6]), .B(a[7]), .ZN(n2927) );
  XOR2_X1 U2524 ( .A(a[4]), .B(n265), .Z(n2939) );
  XNOR2_X1 U2525 ( .A(a[3]), .B(a[4]), .ZN(n2928) );
  XOR2_X1 U2526 ( .A(a[1]), .B(n262), .Z(n2940) );
  XNOR2_X1 U2527 ( .A(a[30]), .B(a[31]), .ZN(n2919) );
  XNOR2_X1 U2528 ( .A(a[0]), .B(a[1]), .ZN(n2929) );
  INV_X1 U2529 ( .A(a[0]), .ZN(n2918) );
  OR2_X1 U2530 ( .A1(n2929), .A2(a[0]), .ZN(n3230) );
  BUF_X1 U2531 ( .A(n351), .Z(n3126) );
  BUF_X1 U2532 ( .A(n348), .Z(n3127) );
  BUF_X1 U2533 ( .A(n354), .Z(n3128) );
  OR2_X1 U2534 ( .A1(n2908), .A2(a[31]), .ZN(n3129) );
  INV_X1 U2535 ( .A(n3129), .ZN(n3130) );
  INV_X1 U2536 ( .A(n3129), .ZN(n3131) );
  XNOR2_X1 U2537 ( .A(n289), .B(a[30]), .ZN(n2908) );
  OR2_X1 U2538 ( .A1(n2931), .A2(n2909), .ZN(n3132) );
  INV_X1 U2539 ( .A(n3132), .ZN(n3133) );
  INV_X1 U2540 ( .A(n3132), .ZN(n3134) );
  XNOR2_X1 U2541 ( .A(n286), .B(a[27]), .ZN(n2909) );
  OR2_X1 U2542 ( .A1(n2932), .A2(n2910), .ZN(n3135) );
  INV_X1 U2543 ( .A(n3135), .ZN(n3136) );
  INV_X1 U2544 ( .A(n3135), .ZN(n3137) );
  XNOR2_X1 U2545 ( .A(n283), .B(a[24]), .ZN(n2910) );
  OR2_X1 U2546 ( .A1(n2933), .A2(n2911), .ZN(n3138) );
  INV_X1 U2547 ( .A(n3138), .ZN(n3139) );
  INV_X1 U2548 ( .A(n3138), .ZN(n3140) );
  OR2_X1 U2549 ( .A1(n2934), .A2(n2912), .ZN(n3141) );
  INV_X1 U2550 ( .A(n3141), .ZN(n3142) );
  INV_X1 U2551 ( .A(n3141), .ZN(n3143) );
  OR2_X1 U2552 ( .A1(n2935), .A2(n2913), .ZN(n3144) );
  INV_X1 U2553 ( .A(n3144), .ZN(n3145) );
  INV_X1 U2554 ( .A(n3144), .ZN(n3146) );
  OR2_X1 U2555 ( .A1(n2936), .A2(n2914), .ZN(n3147) );
  INV_X1 U2556 ( .A(n3147), .ZN(n3148) );
  INV_X1 U2557 ( .A(n3147), .ZN(n3149) );
  OR2_X1 U2558 ( .A1(n2940), .A2(n2918), .ZN(n3150) );
  INV_X1 U2559 ( .A(n3150), .ZN(n3151) );
  INV_X1 U2560 ( .A(n3150), .ZN(n3152) );
  AND2_X1 U2561 ( .A1(n2932), .A2(n3222), .ZN(n3153) );
  INV_X1 U2562 ( .A(n3153), .ZN(n3154) );
  INV_X4 U2563 ( .A(n3153), .ZN(n3155) );
  AND2_X1 U2564 ( .A1(n2931), .A2(n3221), .ZN(n3156) );
  INV_X1 U2565 ( .A(n3156), .ZN(n3157) );
  INV_X4 U2566 ( .A(n3156), .ZN(n3158) );
  AND2_X1 U2567 ( .A1(a[31]), .A2(n3220), .ZN(n3159) );
  INV_X1 U2568 ( .A(n3159), .ZN(n3160) );
  INV_X4 U2569 ( .A(n3159), .ZN(n3161) );
  BUF_X1 U2570 ( .A(n357), .Z(n3162) );
  NAND2_X4 U2571 ( .A1(n2933), .A2(n3223), .ZN(n357) );
  XOR2_X1 U2572 ( .A(n726), .B(n728), .Z(n3163) );
  XOR2_X1 U2573 ( .A(n3163), .B(n523), .Z(product[59]) );
  NAND2_X2 U2574 ( .A1(n726), .A2(n728), .ZN(n3164) );
  NAND2_X1 U2575 ( .A1(n726), .A2(n523), .ZN(n3165) );
  NAND2_X1 U2576 ( .A1(n728), .A2(n523), .ZN(n3166) );
  NAND3_X2 U2577 ( .A1(n3164), .A2(n3165), .A3(n3166), .ZN(n522) );
  XOR2_X1 U2578 ( .A(n725), .B(n722), .Z(n3167) );
  XOR2_X1 U2579 ( .A(n3167), .B(n522), .Z(product[60]) );
  NAND2_X1 U2580 ( .A1(n725), .A2(n722), .ZN(n3168) );
  NAND2_X1 U2581 ( .A1(n725), .A2(n522), .ZN(n3169) );
  NAND2_X1 U2582 ( .A1(n722), .A2(n522), .ZN(n3170) );
  NAND3_X1 U2583 ( .A1(n3168), .A2(n3169), .A3(n3170), .ZN(n521) );
  BUF_X1 U2584 ( .A(n545), .Z(n3171) );
  XOR2_X1 U2585 ( .A(n997), .B(n1014), .Z(n3172) );
  XOR2_X1 U2586 ( .A(n547), .B(n3172), .Z(product[35]) );
  NAND2_X1 U2587 ( .A1(n547), .A2(n997), .ZN(n3173) );
  NAND2_X1 U2588 ( .A1(n547), .A2(n1014), .ZN(n3174) );
  NAND2_X1 U2589 ( .A1(n997), .A2(n1014), .ZN(n3175) );
  NAND3_X2 U2590 ( .A1(n3173), .A2(n3175), .A3(n3174), .ZN(n546) );
  AOI21_X1 U2591 ( .B1(n643), .B2(n706), .A(n640), .ZN(n3176) );
  NAND2_X1 U2592 ( .A1(n651), .A2(n708), .ZN(n3177) );
  INV_X1 U2593 ( .A(n648), .ZN(n3178) );
  AND2_X2 U2594 ( .A1(n3177), .A2(n3178), .ZN(n646) );
  AOI21_X1 U2595 ( .B1(n563), .B2(n686), .A(n560), .ZN(n3179) );
  NAND3_X1 U2596 ( .A1(n3190), .A2(n3192), .A3(n3191), .ZN(n545) );
  AOI21_X2 U2597 ( .B1(n643), .B2(n706), .A(n640), .ZN(n638) );
  OAI21_X1 U2598 ( .B1(n654), .B2(n652), .A(n653), .ZN(n651) );
  INV_X1 U2599 ( .A(n650), .ZN(n648) );
  OAI21_X1 U2600 ( .B1(n644), .B2(n646), .A(n645), .ZN(n643) );
  OAI21_X2 U2601 ( .B1(n566), .B2(n564), .A(n565), .ZN(n563) );
  AOI21_X2 U2602 ( .B1(n563), .B2(n686), .A(n560), .ZN(n558) );
  AOI21_X2 U2603 ( .B1(n587), .B2(n692), .A(n584), .ZN(n582) );
  XOR2_X1 U2604 ( .A(n719), .B(n718), .Z(n3180) );
  XOR2_X1 U2605 ( .A(n520), .B(n3180), .Z(product[62]) );
  NAND2_X1 U2606 ( .A1(n520), .A2(n719), .ZN(n3181) );
  NAND2_X1 U2607 ( .A1(n520), .A2(n718), .ZN(n3182) );
  NAND2_X1 U2608 ( .A1(n719), .A2(n718), .ZN(n3183) );
  NAND3_X1 U2609 ( .A1(n3181), .A2(n3183), .A3(n3182), .ZN(n519) );
  XOR2_X1 U2610 ( .A(n720), .B(n721), .Z(n3184) );
  XOR2_X1 U2611 ( .A(n521), .B(n3184), .Z(product[61]) );
  NAND2_X1 U2612 ( .A1(n521), .A2(n720), .ZN(n3185) );
  NAND2_X1 U2613 ( .A1(n521), .A2(n721), .ZN(n3186) );
  NAND2_X1 U2614 ( .A1(n720), .A2(n721), .ZN(n3187) );
  NAND3_X1 U2615 ( .A1(n3185), .A2(n3187), .A3(n3186), .ZN(n520) );
  BUF_X1 U2616 ( .A(n544), .Z(n3188) );
  XOR2_X1 U2617 ( .A(n996), .B(n979), .Z(n3189) );
  XOR2_X1 U2618 ( .A(n546), .B(n3189), .Z(product[36]) );
  NAND2_X1 U2619 ( .A1(n546), .A2(n996), .ZN(n3190) );
  NAND2_X1 U2620 ( .A1(n546), .A2(n979), .ZN(n3191) );
  NAND2_X1 U2621 ( .A1(n996), .A2(n979), .ZN(n3192) );
  BUF_X1 U2622 ( .A(n635), .Z(n3193) );
  BUF_X1 U2623 ( .A(n627), .Z(n3194) );
  BUF_X1 U2624 ( .A(n579), .Z(n3195) );
  INV_X1 U2625 ( .A(n717), .ZN(n718) );
  NAND3_X1 U2626 ( .A1(n3205), .A2(n3206), .A3(n3207), .ZN(n544) );
  OAI21_X1 U2627 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  AOI21_X2 U2628 ( .B1(n627), .B2(n702), .A(n624), .ZN(n622) );
  XOR2_X1 U2629 ( .A(n582), .B(n494), .Z(product[26]) );
  OAI21_X1 U2630 ( .B1(n582), .B2(n580), .A(n581), .ZN(n579) );
  OAI21_X1 U2631 ( .B1(n630), .B2(n628), .A(n629), .ZN(n627) );
  XOR2_X1 U2632 ( .A(n614), .B(n502), .Z(product[18]) );
  AOI21_X2 U2633 ( .B1(n635), .B2(n704), .A(n632), .ZN(n630) );
  XNOR2_X1 U2634 ( .A(n513), .B(n659), .ZN(product[7]) );
  XOR2_X1 U2635 ( .A(n3179), .B(n488), .Z(product[32]) );
  NOR2_X2 U2636 ( .A1(n2090), .A2(n1373), .ZN(n673) );
  NAND2_X2 U2637 ( .A1(n2090), .A2(n1373), .ZN(n674) );
  OAI21_X1 U2638 ( .B1(n2841), .B2(n345), .A(n2603), .ZN(n2569) );
  XOR2_X1 U2639 ( .A(n2569), .B(n271), .Z(n1988) );
  NOR2_X2 U2640 ( .A1(n1339), .A2(n1344), .ZN(n641) );
  XOR2_X1 U2641 ( .A(n773), .B(n782), .Z(n3196) );
  XOR2_X1 U2642 ( .A(n3196), .B(n531), .Z(product[51]) );
  NAND2_X2 U2643 ( .A1(n773), .A2(n782), .ZN(n3197) );
  NAND2_X1 U2644 ( .A1(n773), .A2(n531), .ZN(n3198) );
  NAND2_X1 U2645 ( .A1(n782), .A2(n531), .ZN(n3199) );
  NAND3_X2 U2646 ( .A1(n3197), .A2(n3198), .A3(n3199), .ZN(n530) );
  XOR2_X1 U2647 ( .A(n765), .B(n772), .Z(n3200) );
  XOR2_X1 U2648 ( .A(n3200), .B(n530), .Z(product[52]) );
  NAND2_X1 U2649 ( .A1(n765), .A2(n772), .ZN(n3201) );
  NAND2_X1 U2650 ( .A1(n765), .A2(n530), .ZN(n3202) );
  NAND2_X1 U2651 ( .A1(n772), .A2(n530), .ZN(n3203) );
  NAND3_X1 U2652 ( .A1(n3201), .A2(n3202), .A3(n3203), .ZN(n529) );
  XOR2_X1 U2653 ( .A(n961), .B(n978), .Z(n3204) );
  XOR2_X1 U2654 ( .A(n3204), .B(n3171), .Z(product[37]) );
  NAND2_X2 U2655 ( .A1(n961), .A2(n978), .ZN(n3205) );
  NAND2_X1 U2656 ( .A1(n961), .A2(n545), .ZN(n3206) );
  NAND2_X1 U2657 ( .A1(n978), .A2(n545), .ZN(n3207) );
  XOR2_X1 U2658 ( .A(n944), .B(n960), .Z(n3208) );
  XOR2_X1 U2659 ( .A(n3208), .B(n3188), .Z(product[38]) );
  NAND2_X1 U2660 ( .A1(n944), .A2(n960), .ZN(n3209) );
  NAND2_X1 U2661 ( .A1(n944), .A2(n544), .ZN(n3210) );
  NAND2_X1 U2662 ( .A1(n960), .A2(n544), .ZN(n3211) );
  NAND3_X1 U2663 ( .A1(n3209), .A2(n3210), .A3(n3211), .ZN(n543) );
  AOI21_X1 U2664 ( .B1(n555), .B2(n684), .A(n552), .ZN(n3212) );
  OR2_X1 U2665 ( .A1(n2841), .A2(n342), .ZN(n3213) );
  NAND2_X1 U2666 ( .A1(n3213), .A2(n2671), .ZN(n2637) );
  BUF_X1 U2667 ( .A(n595), .Z(n3214) );
  INV_X8 U2668 ( .A(n390), .ZN(n2841) );
  INV_X1 U2669 ( .A(n1400), .ZN(n2671) );
  XNOR2_X1 U2670 ( .A(n3193), .B(n507), .ZN(product[13]) );
  XOR2_X1 U2671 ( .A(n630), .B(n506), .Z(product[14]) );
  NAND2_X4 U2672 ( .A1(n2934), .A2(n3224), .ZN(n354) );
  XOR2_X1 U2673 ( .A(n3176), .B(n508), .Z(product[12]) );
  XOR2_X1 U2674 ( .A(n2365), .B(n280), .Z(n1883) );
  OR2_X4 U2675 ( .A1(n2928), .A2(n3229), .ZN(n3231) );
  INV_X8 U2676 ( .A(n3231), .ZN(n315) );
  AOI21_X4 U2677 ( .B1(n603), .B2(n696), .A(n600), .ZN(n598) );
  INV_X1 U2678 ( .A(n649), .ZN(n708) );
  XOR2_X1 U2679 ( .A(n2637), .B(n268), .Z(n2023) );
  NOR2_X1 U2680 ( .A1(n1351), .A2(n1356), .ZN(n649) );
  NAND2_X2 U2681 ( .A1(n1351), .A2(n1356), .ZN(n650) );
  OR2_X4 U2682 ( .A1(n2927), .A2(n3228), .ZN(n3232) );
  INV_X8 U2683 ( .A(n3232), .ZN(n317) );
  OR2_X4 U2684 ( .A1(n2937), .A2(n2915), .ZN(n3215) );
  INV_X32 U2685 ( .A(n3215), .ZN(n297) );
  AOI22_X1 U2686 ( .A1(n295), .A2(n393), .B1(n317), .B2(n390), .ZN(n2670) );
  OAI21_X1 U2687 ( .B1(n2840), .B2(n342), .A(n2670), .ZN(n2636) );
  XOR2_X1 U2688 ( .A(n2636), .B(n268), .Z(n2022) );
  INV_X2 U2689 ( .A(n293), .ZN(n3216) );
  INV_X8 U2690 ( .A(n3216), .ZN(n3217) );
  NOR2_X2 U2691 ( .A1(n2939), .A2(n2917), .ZN(n293) );
  XNOR2_X1 U2692 ( .A(n3214), .B(n497), .ZN(product[23]) );
  XNOR2_X1 U2693 ( .A(n603), .B(n499), .ZN(product[21]) );
  OAI21_X2 U2694 ( .B1(n660), .B2(n662), .A(n661), .ZN(n659) );
  NOR2_X2 U2695 ( .A1(n1365), .A2(n2087), .ZN(n660) );
  OAI21_X1 U2696 ( .B1(n2841), .B2(n339), .A(n2739), .ZN(n2705) );
  INV_X1 U2697 ( .A(n1403), .ZN(n2739) );
  OAI21_X2 U2698 ( .B1(n606), .B2(n604), .A(n605), .ZN(n603) );
  XOR2_X1 U2699 ( .A(n598), .B(n498), .Z(product[22]) );
  OAI21_X2 U2700 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  NAND2_X4 U2701 ( .A1(n2935), .A2(n3225), .ZN(n351) );
  OR2_X4 U2702 ( .A1(n2938), .A2(n2916), .ZN(n3218) );
  INV_X32 U2703 ( .A(n3218), .ZN(n295) );
  XNOR2_X1 U2704 ( .A(n519), .B(n3219), .ZN(product[63]) );
  INV_X32 U2705 ( .A(n485), .ZN(n3219) );
  XNOR2_X1 U2706 ( .A(n611), .B(n501), .ZN(product[19]) );
  NAND2_X4 U2707 ( .A1(n2940), .A2(a[0]), .ZN(n336) );
  OAI21_X2 U2708 ( .B1(n614), .B2(n612), .A(n613), .ZN(n611) );
  OAI21_X1 U2709 ( .B1(n574), .B2(n572), .A(n573), .ZN(n571) );
  NAND2_X4 U2710 ( .A1(n2936), .A2(n3226), .ZN(n348) );
  XNOR2_X1 U2711 ( .A(n563), .B(n489), .ZN(product[31]) );
  XNOR2_X1 U2712 ( .A(n619), .B(n503), .ZN(product[17]) );
  NAND2_X1 U2713 ( .A1(n715), .A2(n682), .ZN(n518) );
  XOR2_X1 U2714 ( .A(n566), .B(n490), .Z(product[30]) );
  XOR2_X1 U2715 ( .A(n622), .B(n504), .Z(product[16]) );
  NOR2_X1 U2716 ( .A1(n2093), .A2(n262), .ZN(n681) );
  AOI21_X2 U2717 ( .B1(n571), .B2(n688), .A(n568), .ZN(n566) );
  AOI21_X2 U2718 ( .B1(n579), .B2(n690), .A(n576), .ZN(n574) );
  OAI21_X2 U2719 ( .B1(n622), .B2(n620), .A(n621), .ZN(n619) );
  XNOR2_X1 U2720 ( .A(n571), .B(n491), .ZN(product[29]) );
  XNOR2_X1 U2721 ( .A(n651), .B(n511), .ZN(product[9]) );
  XNOR2_X1 U2722 ( .A(n643), .B(n509), .ZN(product[11]) );
  XOR2_X1 U2723 ( .A(n3212), .B(n486), .Z(product[34]) );
  OAI21_X1 U2724 ( .B1(n2841), .B2(n336), .A(n2807), .ZN(n2773) );
  XOR2_X1 U2725 ( .A(n2773), .B(n262), .Z(n2093) );
  NAND2_X2 U2726 ( .A1(n2093), .A2(n262), .ZN(n682) );
  NAND2_X4 U2727 ( .A1(n2937), .A2(n3227), .ZN(n345) );
  NAND2_X4 U2728 ( .A1(n2938), .A2(n3228), .ZN(n342) );
  XNOR2_X1 U2729 ( .A(n3195), .B(n493), .ZN(product[27]) );
  XNOR2_X1 U2730 ( .A(n3194), .B(n505), .ZN(product[15]) );
  XNOR2_X1 U2731 ( .A(n555), .B(n487), .ZN(product[33]) );
  XNOR2_X1 U2732 ( .A(n587), .B(n495), .ZN(product[25]) );
  XOR2_X1 U2733 ( .A(n574), .B(n492), .Z(product[28]) );
  XOR2_X1 U2734 ( .A(n510), .B(n646), .Z(product[10]) );
  AOI21_X2 U2735 ( .B1(n555), .B2(n684), .A(n552), .ZN(n550) );
  NAND2_X4 U2736 ( .A1(n2939), .A2(n3229), .ZN(n339) );
  OAI21_X1 U2737 ( .B1(n550), .B2(n548), .A(n549), .ZN(n547) );
  OAI21_X2 U2738 ( .B1(n558), .B2(n556), .A(n557), .ZN(n555) );
  OAI21_X2 U2739 ( .B1(n590), .B2(n588), .A(n589), .ZN(n587) );
  INV_X2 U2740 ( .A(n518), .ZN(product[0]) );
  INV_X2 U2741 ( .A(n941), .ZN(n959) );
  INV_X2 U2742 ( .A(n907), .ZN(n908) );
  INV_X2 U2743 ( .A(n891), .ZN(n892) );
  INV_X2 U2744 ( .A(n848), .ZN(n862) );
  INV_X2 U2745 ( .A(n811), .ZN(n823) );
  INV_X2 U2746 ( .A(n780), .ZN(n790) );
  INV_X2 U2747 ( .A(n755), .ZN(n763) );
  INV_X2 U2748 ( .A(n736), .ZN(n742) );
  INV_X2 U2749 ( .A(n723), .ZN(n727) );
  INV_X2 U2750 ( .A(n1720), .ZN(n716) );
  INV_X2 U2751 ( .A(n681), .ZN(n715) );
  INV_X2 U2752 ( .A(n668), .ZN(n713) );
  INV_X2 U2753 ( .A(n660), .ZN(n711) );
  INV_X2 U2754 ( .A(n652), .ZN(n709) );
  INV_X2 U2755 ( .A(n644), .ZN(n707) );
  INV_X2 U2756 ( .A(n636), .ZN(n705) );
  INV_X2 U2757 ( .A(n628), .ZN(n703) );
  INV_X2 U2758 ( .A(n620), .ZN(n701) );
  INV_X2 U2759 ( .A(n612), .ZN(n699) );
  INV_X2 U2760 ( .A(n604), .ZN(n697) );
  INV_X2 U2761 ( .A(n596), .ZN(n695) );
  INV_X2 U2762 ( .A(n588), .ZN(n693) );
  INV_X2 U2763 ( .A(n580), .ZN(n691) );
  INV_X2 U2764 ( .A(n572), .ZN(n689) );
  INV_X2 U2765 ( .A(n564), .ZN(n687) );
  INV_X2 U2766 ( .A(n556), .ZN(n685) );
  INV_X2 U2767 ( .A(n548), .ZN(n683) );
  INV_X2 U2768 ( .A(n682), .ZN(n680) );
  INV_X2 U2769 ( .A(n678), .ZN(n679) );
  INV_X2 U2770 ( .A(n2091), .ZN(n676) );
  INV_X2 U2771 ( .A(n674), .ZN(n672) );
  INV_X2 U2772 ( .A(n673), .ZN(n714) );
  INV_X2 U2773 ( .A(n666), .ZN(n664) );
  INV_X2 U2774 ( .A(n665), .ZN(n712) );
  INV_X2 U2775 ( .A(n658), .ZN(n656) );
  INV_X2 U2776 ( .A(n657), .ZN(n710) );
  INV_X2 U2777 ( .A(n642), .ZN(n640) );
  INV_X2 U2778 ( .A(n641), .ZN(n706) );
  INV_X2 U2779 ( .A(n634), .ZN(n632) );
  INV_X2 U2780 ( .A(n633), .ZN(n704) );
  INV_X2 U2781 ( .A(n626), .ZN(n624) );
  INV_X2 U2782 ( .A(n625), .ZN(n702) );
  INV_X2 U2783 ( .A(n618), .ZN(n616) );
  INV_X2 U2784 ( .A(n617), .ZN(n700) );
  INV_X2 U2785 ( .A(n610), .ZN(n608) );
  INV_X2 U2786 ( .A(n609), .ZN(n698) );
  INV_X2 U2787 ( .A(n602), .ZN(n600) );
  INV_X2 U2788 ( .A(n601), .ZN(n696) );
  INV_X2 U2789 ( .A(n594), .ZN(n592) );
  INV_X2 U2790 ( .A(n593), .ZN(n694) );
  INV_X2 U2791 ( .A(n586), .ZN(n584) );
  INV_X2 U2792 ( .A(n585), .ZN(n692) );
  INV_X2 U2793 ( .A(n578), .ZN(n576) );
  INV_X2 U2794 ( .A(n577), .ZN(n690) );
  INV_X2 U2795 ( .A(n570), .ZN(n568) );
  INV_X2 U2796 ( .A(n569), .ZN(n688) );
  INV_X2 U2797 ( .A(n562), .ZN(n560) );
  INV_X2 U2798 ( .A(n561), .ZN(n686) );
  INV_X2 U2799 ( .A(n554), .ZN(n552) );
  INV_X2 U2800 ( .A(n553), .ZN(n684) );
  INV_X2 U2801 ( .A(n2873), .ZN(n2839) );
  INV_X2 U2802 ( .A(n2872), .ZN(n2838) );
  INV_X2 U2803 ( .A(n2871), .ZN(n2837) );
  INV_X2 U2804 ( .A(n2870), .ZN(n2836) );
  INV_X2 U2805 ( .A(n2869), .ZN(n2835) );
  INV_X2 U2806 ( .A(n2868), .ZN(n2834) );
  INV_X2 U2807 ( .A(n2867), .ZN(n2833) );
  INV_X2 U2808 ( .A(n2866), .ZN(n2832) );
  INV_X2 U2809 ( .A(n2865), .ZN(n2831) );
  INV_X2 U2810 ( .A(n2864), .ZN(n2830) );
  INV_X2 U2811 ( .A(n2863), .ZN(n2829) );
  INV_X2 U2812 ( .A(n2862), .ZN(n2828) );
  INV_X2 U2813 ( .A(n2861), .ZN(n2827) );
  INV_X2 U2814 ( .A(n2860), .ZN(n2826) );
  INV_X2 U2815 ( .A(n2859), .ZN(n2825) );
  INV_X2 U2816 ( .A(n2858), .ZN(n2824) );
  INV_X2 U2817 ( .A(n2857), .ZN(n2823) );
  INV_X2 U2818 ( .A(n2856), .ZN(n2822) );
  INV_X2 U2819 ( .A(n2855), .ZN(n2821) );
  INV_X2 U2820 ( .A(n2854), .ZN(n2820) );
  INV_X2 U2821 ( .A(n2853), .ZN(n2819) );
  INV_X2 U2822 ( .A(n2852), .ZN(n2818) );
  INV_X2 U2823 ( .A(n2851), .ZN(n2817) );
  INV_X2 U2824 ( .A(n2850), .ZN(n2816) );
  INV_X2 U2825 ( .A(n2849), .ZN(n2815) );
  INV_X2 U2826 ( .A(n2848), .ZN(n2814) );
  INV_X2 U2827 ( .A(n2847), .ZN(n2813) );
  INV_X2 U2828 ( .A(n2846), .ZN(n2812) );
  INV_X2 U2829 ( .A(n2845), .ZN(n2811) );
  INV_X2 U2830 ( .A(n2844), .ZN(n2810) );
  INV_X2 U2831 ( .A(n2843), .ZN(n2809) );
  INV_X2 U2832 ( .A(n1406), .ZN(n2807) );
  AOI22_X2 U2833 ( .A1(n3152), .A2(n393), .B1(n313), .B2(n390), .ZN(n2806) );
  INV_X2 U2834 ( .A(n3230), .ZN(n313) );
  AOI22_X2 U2835 ( .A1(n3217), .A2(n393), .B1(n315), .B2(n390), .ZN(n2738) );
  INV_X2 U2836 ( .A(n2917), .ZN(n3229) );
  INV_X2 U2837 ( .A(n2916), .ZN(n3228) );
  INV_X2 U2838 ( .A(n1397), .ZN(n2603) );
  AOI22_X2 U2839 ( .A1(n297), .A2(n393), .B1(n319), .B2(n390), .ZN(n2602) );
  INV_X2 U2840 ( .A(n3233), .ZN(n319) );
  OR2_X2 U2841 ( .A1(n2926), .A2(n3227), .ZN(n3233) );
  INV_X2 U2842 ( .A(n2915), .ZN(n3227) );
  INV_X2 U2843 ( .A(n1394), .ZN(n2535) );
  AOI22_X2 U2844 ( .A1(n3149), .A2(n393), .B1(n321), .B2(n390), .ZN(n2534) );
  INV_X2 U2845 ( .A(n3234), .ZN(n321) );
  OR2_X2 U2846 ( .A1(n2925), .A2(n3226), .ZN(n3234) );
  INV_X2 U2847 ( .A(n2914), .ZN(n3226) );
  INV_X2 U2848 ( .A(n1391), .ZN(n2467) );
  AOI22_X2 U2849 ( .A1(n3146), .A2(n393), .B1(n323), .B2(n390), .ZN(n2466) );
  INV_X2 U2850 ( .A(n3235), .ZN(n323) );
  OR2_X2 U2851 ( .A1(n2924), .A2(n3225), .ZN(n3235) );
  INV_X2 U2852 ( .A(n2913), .ZN(n3225) );
  INV_X2 U2853 ( .A(n1388), .ZN(n2399) );
  AOI22_X2 U2854 ( .A1(n3143), .A2(n393), .B1(n325), .B2(n390), .ZN(n2398) );
  INV_X2 U2855 ( .A(n3236), .ZN(n325) );
  OR2_X2 U2856 ( .A1(n2923), .A2(n3224), .ZN(n3236) );
  INV_X2 U2857 ( .A(n2912), .ZN(n3224) );
  INV_X2 U2858 ( .A(n1385), .ZN(n2331) );
  AOI22_X2 U2859 ( .A1(n3140), .A2(n393), .B1(n327), .B2(n390), .ZN(n2330) );
  INV_X2 U2860 ( .A(n3237), .ZN(n327) );
  OR2_X2 U2861 ( .A1(n2922), .A2(n3223), .ZN(n3237) );
  INV_X2 U2862 ( .A(n2911), .ZN(n3223) );
  INV_X2 U2863 ( .A(n1382), .ZN(n2263) );
  AOI22_X2 U2864 ( .A1(n3137), .A2(n393), .B1(n329), .B2(n390), .ZN(n2262) );
  INV_X2 U2865 ( .A(n3238), .ZN(n329) );
  OR2_X2 U2866 ( .A1(n2921), .A2(n3222), .ZN(n3238) );
  INV_X2 U2867 ( .A(n2910), .ZN(n3222) );
  INV_X2 U2868 ( .A(n1379), .ZN(n2195) );
  AOI22_X2 U2869 ( .A1(n3134), .A2(n393), .B1(n331), .B2(n390), .ZN(n2194) );
  INV_X2 U2870 ( .A(n3239), .ZN(n331) );
  OR2_X2 U2871 ( .A1(n2920), .A2(n3221), .ZN(n3239) );
  INV_X2 U2872 ( .A(n2909), .ZN(n3221) );
  INV_X2 U2873 ( .A(n1376), .ZN(n2127) );
  AOI22_X2 U2874 ( .A1(n3130), .A2(n393), .B1(n333), .B2(n390), .ZN(n2126) );
  INV_X2 U2875 ( .A(n3240), .ZN(n333) );
  OR2_X2 U2876 ( .A1(n2919), .A2(n3220), .ZN(n3240) );
  INV_X2 U2877 ( .A(n2908), .ZN(n3220) );
  INV_X2 U2878 ( .A(n262), .ZN(n2059) );
  INV_X2 U2879 ( .A(n265), .ZN(n2024) );
  INV_X2 U2880 ( .A(n268), .ZN(n1989) );
  INV_X2 U2881 ( .A(n271), .ZN(n1954) );
  INV_X2 U2882 ( .A(n274), .ZN(n1919) );
  INV_X2 U2883 ( .A(n277), .ZN(n1884) );
  INV_X2 U2884 ( .A(n280), .ZN(n1849) );
  INV_X2 U2885 ( .A(n283), .ZN(n1814) );
  INV_X2 U2886 ( .A(n286), .ZN(n1779) );
  INV_X2 U2887 ( .A(n289), .ZN(n1745) );
  INV_X2 U2888 ( .A(n1686), .ZN(n1719) );
  INV_X2 U2889 ( .A(n1682), .ZN(n1718) );
  INV_X2 U2890 ( .A(n1679), .ZN(n1717) );
  INV_X2 U2891 ( .A(n1668), .ZN(n1715) );
  INV_X2 U2892 ( .A(n1663), .ZN(n1714) );
  INV_X2 U2893 ( .A(n1660), .ZN(n1713) );
  INV_X2 U2894 ( .A(n1652), .ZN(n1712) );
  INV_X2 U2895 ( .A(n1649), .ZN(n1711) );
  INV_X2 U2896 ( .A(n1637), .ZN(n1709) );
  INV_X2 U2897 ( .A(n1621), .ZN(n1707) );
  INV_X2 U2898 ( .A(n1607), .ZN(n1705) );
  INV_X2 U2899 ( .A(n1592), .ZN(n1703) );
  INV_X2 U2900 ( .A(n1581), .ZN(n1702) );
  INV_X2 U2901 ( .A(n1576), .ZN(n1701) );
  INV_X2 U2902 ( .A(n1561), .ZN(n1700) );
  INV_X2 U2903 ( .A(n1556), .ZN(n1699) );
  INV_X2 U2904 ( .A(n1543), .ZN(n1698) );
  INV_X2 U2905 ( .A(n1538), .ZN(n1697) );
  INV_X2 U2906 ( .A(n1523), .ZN(n1696) );
  INV_X2 U2907 ( .A(n1518), .ZN(n1695) );
  INV_X2 U2908 ( .A(n1496), .ZN(n1693) );
  INV_X2 U2909 ( .A(n1474), .ZN(n1691) );
  INV_X2 U2910 ( .A(n1459), .ZN(n1690) );
  INV_X2 U2911 ( .A(n1450), .ZN(n1689) );
  INV_X2 U2912 ( .A(n1684), .ZN(n1685) );
  INV_X2 U2913 ( .A(n1676), .ZN(n1675) );
  INV_X2 U2914 ( .A(n1674), .ZN(n1672) );
  INV_X2 U2915 ( .A(n1673), .ZN(n1716) );
  INV_X2 U2916 ( .A(n1655), .ZN(n1654) );
  INV_X2 U2917 ( .A(n1648), .ZN(n1646) );
  INV_X2 U2918 ( .A(n1647), .ZN(n1645) );
  INV_X2 U2919 ( .A(n1643), .ZN(n1641) );
  INV_X2 U2920 ( .A(n1642), .ZN(n1710) );
  INV_X2 U2921 ( .A(n1630), .ZN(n1632) );
  INV_X2 U2922 ( .A(n1629), .ZN(n1631) );
  INV_X2 U2923 ( .A(n1627), .ZN(n1625) );
  INV_X2 U2924 ( .A(n1626), .ZN(n1708) );
  INV_X2 U2925 ( .A(n1613), .ZN(n1611) );
  INV_X2 U2926 ( .A(n1612), .ZN(n1706) );
  INV_X2 U2927 ( .A(n1600), .ZN(n1599) );
  INV_X2 U2928 ( .A(n1598), .ZN(n1596) );
  INV_X2 U2929 ( .A(n1597), .ZN(n1704) );
  INV_X2 U2930 ( .A(n1587), .ZN(n1589) );
  INV_X2 U2931 ( .A(n1586), .ZN(n1588) );
  INV_X2 U2932 ( .A(n1569), .ZN(n1571) );
  INV_X2 U2933 ( .A(n1568), .ZN(n1570) );
  INV_X2 U2934 ( .A(n1551), .ZN(n1549) );
  INV_X2 U2935 ( .A(n1550), .ZN(n1548) );
  INV_X2 U2936 ( .A(n1529), .ZN(n1531) );
  INV_X2 U2937 ( .A(n1528), .ZN(n1530) );
  INV_X2 U2938 ( .A(n1513), .ZN(n1511) );
  INV_X2 U2939 ( .A(n1512), .ZN(n1510) );
  INV_X2 U2940 ( .A(n1506), .ZN(n1504) );
  INV_X2 U2941 ( .A(n1505), .ZN(n1694) );
  INV_X2 U2942 ( .A(n1489), .ZN(n1491) );
  INV_X2 U2943 ( .A(n1488), .ZN(n1490) );
  INV_X2 U2944 ( .A(n1484), .ZN(n1482) );
  INV_X2 U2945 ( .A(n1483), .ZN(n1692) );
  INV_X2 U2946 ( .A(n1469), .ZN(n1471) );
  INV_X2 U2947 ( .A(n1468), .ZN(n1470) );
  INV_X2 U2948 ( .A(n484), .ZN(n1440) );
endmodule


module mul32_2_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n262, n265, n268, n271, n274, n277, n280, n283, n286, n289, n293,
         n295, n297, n299, n313, n315, n317, n319, n321, n323, n325, n327,
         n329, n331, n333, n336, n339, n342, n345, n348, n351, n354, n357,
         n360, n368, n370, n374, n376, n378, n380, n382, n384, n386, n388,
         n390, n393, n397, n400, n403, n406, n409, n412, n415, n418, n421,
         n424, n427, n430, n433, n436, n439, n442, n445, n448, n451, n454,
         n457, n460, n463, n466, n469, n472, n475, n478, n481, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n552,
         n553, n554, n555, n556, n557, n558, n560, n561, n562, n563, n564,
         n565, n566, n568, n569, n570, n571, n572, n573, n574, n576, n577,
         n578, n579, n580, n581, n582, n584, n585, n586, n587, n588, n589,
         n590, n592, n593, n594, n595, n596, n597, n598, n600, n601, n602,
         n603, n604, n605, n606, n608, n609, n610, n611, n612, n613, n614,
         n616, n617, n618, n619, n620, n621, n622, n624, n625, n626, n627,
         n628, n629, n630, n632, n633, n634, n635, n636, n637, n638, n640,
         n641, n642, n643, n644, n645, n646, n648, n649, n650, n651, n652,
         n653, n654, n656, n657, n658, n659, n660, n661, n662, n664, n665,
         n666, n667, n668, n669, n670, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1376, n1377, n1379, n1380, n1382, n1383, n1385, n1386, n1388,
         n1389, n1391, n1392, n1394, n1395, n1397, n1398, n1400, n1401, n1403,
         n1404, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1518, n1519,
         n1520, n1521, n1522, n1523, n1526, n1527, n1528, n1529, n1530, n1531,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1564, n1565, n1568, n1569, n1570, n1571,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1584, n1585,
         n1586, n1587, n1588, n1589, n1592, n1593, n1594, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1620, n1621,
         n1622, n1623, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1635, n1636, n1637, n1638, n1639, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248;
  assign n262 = a[2];
  assign n265 = a[5];
  assign n268 = a[8];
  assign n271 = a[11];
  assign n274 = a[14];
  assign n277 = a[17];
  assign n280 = a[20];
  assign n283 = a[23];
  assign n286 = a[26];
  assign n289 = a[29];
  assign n390 = b[0];
  assign n393 = b[1];
  assign n397 = b[2];
  assign n400 = b[3];
  assign n403 = b[4];
  assign n406 = b[5];
  assign n409 = b[6];
  assign n412 = b[7];
  assign n415 = b[8];
  assign n418 = b[9];
  assign n421 = b[10];
  assign n424 = b[11];
  assign n427 = b[12];
  assign n430 = b[13];
  assign n433 = b[14];
  assign n436 = b[15];
  assign n439 = b[16];
  assign n442 = b[17];
  assign n445 = b[18];
  assign n448 = b[19];
  assign n451 = b[20];
  assign n454 = b[21];
  assign n457 = b[22];
  assign n460 = b[23];
  assign n463 = b[24];
  assign n466 = b[25];
  assign n469 = b[26];
  assign n472 = b[27];
  assign n475 = b[28];
  assign n478 = b[29];
  assign n481 = b[30];
  assign n484 = b[31];

  XOR2_X2 U304 ( .A(n717), .B(n716), .Z(n485) );
  FA_X1 U306 ( .A(n720), .B(n721), .CI(n521), .CO(n520), .S(product[61]) );
  FA_X1 U307 ( .A(n725), .B(n722), .CI(n522), .CO(n521), .S(product[60]) );
  FA_X1 U308 ( .A(n726), .B(n728), .CI(n523), .CO(n522), .S(product[59]) );
  FA_X1 U314 ( .A(n744), .B(n749), .CI(n527), .CO(n526), .S(product[55]) );
  FA_X1 U315 ( .A(n750), .B(n757), .CI(n528), .CO(n527), .S(product[54]) );
  FA_X1 U316 ( .A(n758), .B(n764), .CI(n529), .CO(n528), .S(product[53]) );
  FA_X1 U317 ( .A(n765), .B(n772), .CI(n530), .CO(n529), .S(product[52]) );
  FA_X1 U318 ( .A(n773), .B(n782), .CI(n531), .CO(n530), .S(product[51]) );
  FA_X1 U319 ( .A(n783), .B(n791), .CI(n532), .CO(n531), .S(product[50]) );
  FA_X1 U320 ( .A(n792), .B(n801), .CI(n533), .CO(n532), .S(product[49]) );
  FA_X1 U324 ( .A(n837), .B(n850), .CI(n537), .CO(n536), .S(product[45]) );
  FA_X1 U325 ( .A(n851), .B(n863), .CI(n538), .CO(n537), .S(product[44]) );
  FA_X1 U326 ( .A(n864), .B(n877), .CI(n539), .CO(n538), .S(product[43]) );
  FA_X1 U327 ( .A(n878), .B(n893), .CI(n540), .CO(n539), .S(product[42]) );
  FA_X1 U328 ( .A(n894), .B(n909), .CI(n541), .CO(n540), .S(product[41]) );
  FA_X1 U329 ( .A(n910), .B(n925), .CI(n542), .CO(n541), .S(product[40]) );
  FA_X1 U330 ( .A(n926), .B(n943), .CI(n543), .CO(n542), .S(product[39]) );
  FA_X1 U334 ( .A(n997), .B(n1014), .CI(n547), .CO(n546), .S(product[35]) );
  NAND2_X4 U337 ( .A1(n683), .A2(n549), .ZN(n486) );
  NOR2_X4 U339 ( .A1(n1015), .A2(n1032), .ZN(n548) );
  NAND2_X4 U340 ( .A1(n1015), .A2(n1032), .ZN(n549) );
  NAND2_X4 U345 ( .A1(n684), .A2(n554), .ZN(n487) );
  NOR2_X4 U347 ( .A1(n1033), .A2(n1050), .ZN(n553) );
  NAND2_X4 U348 ( .A1(n1033), .A2(n1050), .ZN(n554) );
  XOR2_X2 U349 ( .A(n558), .B(n488), .Z(product[32]) );
  NAND2_X4 U351 ( .A1(n685), .A2(n557), .ZN(n488) );
  NOR2_X4 U353 ( .A1(n1051), .A2(n1068), .ZN(n556) );
  NAND2_X4 U354 ( .A1(n1051), .A2(n1068), .ZN(n557) );
  AOI21_X4 U356 ( .B1(n563), .B2(n686), .A(n560), .ZN(n558) );
  NAND2_X4 U359 ( .A1(n686), .A2(n562), .ZN(n489) );
  NOR2_X4 U361 ( .A1(n1069), .A2(n1086), .ZN(n561) );
  NAND2_X4 U362 ( .A1(n1069), .A2(n1086), .ZN(n562) );
  NAND2_X4 U365 ( .A1(n687), .A2(n565), .ZN(n490) );
  NOR2_X4 U367 ( .A1(n1087), .A2(n1104), .ZN(n564) );
  NAND2_X4 U368 ( .A1(n1087), .A2(n1104), .ZN(n565) );
  NAND2_X4 U373 ( .A1(n688), .A2(n570), .ZN(n491) );
  NOR2_X4 U375 ( .A1(n1105), .A2(n1122), .ZN(n569) );
  NAND2_X4 U376 ( .A1(n1105), .A2(n1122), .ZN(n570) );
  XOR2_X2 U377 ( .A(n574), .B(n492), .Z(product[28]) );
  NAND2_X4 U379 ( .A1(n689), .A2(n573), .ZN(n492) );
  NOR2_X4 U381 ( .A1(n1123), .A2(n1140), .ZN(n572) );
  NAND2_X4 U382 ( .A1(n1123), .A2(n1140), .ZN(n573) );
  AOI21_X4 U384 ( .B1(n579), .B2(n690), .A(n576), .ZN(n574) );
  NAND2_X4 U387 ( .A1(n690), .A2(n578), .ZN(n493) );
  NOR2_X4 U389 ( .A1(n1141), .A2(n1158), .ZN(n577) );
  NAND2_X4 U390 ( .A1(n1141), .A2(n1158), .ZN(n578) );
  XOR2_X2 U391 ( .A(n582), .B(n494), .Z(product[26]) );
  NAND2_X4 U393 ( .A1(n691), .A2(n581), .ZN(n494) );
  NOR2_X4 U395 ( .A1(n1159), .A2(n1174), .ZN(n580) );
  NAND2_X4 U396 ( .A1(n1159), .A2(n1174), .ZN(n581) );
  XNOR2_X2 U397 ( .A(n587), .B(n495), .ZN(product[25]) );
  AOI21_X4 U398 ( .B1(n587), .B2(n692), .A(n584), .ZN(n582) );
  NAND2_X4 U401 ( .A1(n692), .A2(n586), .ZN(n495) );
  NOR2_X4 U403 ( .A1(n1175), .A2(n1190), .ZN(n585) );
  NAND2_X4 U404 ( .A1(n1175), .A2(n1190), .ZN(n586) );
  XOR2_X2 U405 ( .A(n590), .B(n496), .Z(product[24]) );
  OAI21_X4 U406 ( .B1(n590), .B2(n588), .A(n589), .ZN(n587) );
  NAND2_X4 U407 ( .A1(n693), .A2(n589), .ZN(n496) );
  NOR2_X4 U409 ( .A1(n1191), .A2(n1206), .ZN(n588) );
  NAND2_X4 U412 ( .A1(n1191), .A2(n1206), .ZN(n589) );
  XNOR2_X2 U413 ( .A(n595), .B(n497), .ZN(product[23]) );
  AOI21_X4 U414 ( .B1(n595), .B2(n694), .A(n592), .ZN(n590) );
  NAND2_X4 U417 ( .A1(n694), .A2(n594), .ZN(n497) );
  NOR2_X4 U419 ( .A1(n1207), .A2(n1220), .ZN(n593) );
  NAND2_X4 U420 ( .A1(n1207), .A2(n1220), .ZN(n594) );
  XOR2_X2 U421 ( .A(n598), .B(n498), .Z(product[22]) );
  OAI21_X4 U422 ( .B1(n598), .B2(n596), .A(n597), .ZN(n595) );
  NAND2_X4 U423 ( .A1(n695), .A2(n597), .ZN(n498) );
  NOR2_X4 U425 ( .A1(n1221), .A2(n1234), .ZN(n596) );
  NAND2_X4 U426 ( .A1(n1221), .A2(n1234), .ZN(n597) );
  XNOR2_X2 U427 ( .A(n603), .B(n499), .ZN(product[21]) );
  AOI21_X4 U428 ( .B1(n603), .B2(n696), .A(n600), .ZN(n598) );
  NAND2_X4 U431 ( .A1(n696), .A2(n602), .ZN(n499) );
  NOR2_X4 U433 ( .A1(n1235), .A2(n1248), .ZN(n601) );
  NAND2_X4 U434 ( .A1(n1235), .A2(n1248), .ZN(n602) );
  XOR2_X2 U435 ( .A(n606), .B(n500), .Z(product[20]) );
  OAI21_X4 U436 ( .B1(n606), .B2(n604), .A(n605), .ZN(n603) );
  NAND2_X4 U437 ( .A1(n697), .A2(n605), .ZN(n500) );
  NOR2_X4 U439 ( .A1(n1249), .A2(n1260), .ZN(n604) );
  NAND2_X4 U440 ( .A1(n1249), .A2(n1260), .ZN(n605) );
  AOI21_X4 U442 ( .B1(n611), .B2(n698), .A(n608), .ZN(n606) );
  NAND2_X4 U445 ( .A1(n698), .A2(n610), .ZN(n501) );
  NOR2_X4 U447 ( .A1(n1261), .A2(n1272), .ZN(n609) );
  NAND2_X4 U448 ( .A1(n1261), .A2(n1272), .ZN(n610) );
  XOR2_X2 U449 ( .A(n614), .B(n502), .Z(product[18]) );
  NAND2_X4 U451 ( .A1(n699), .A2(n613), .ZN(n502) );
  NOR2_X4 U453 ( .A1(n1273), .A2(n1284), .ZN(n612) );
  NAND2_X4 U454 ( .A1(n1273), .A2(n1284), .ZN(n613) );
  AOI21_X4 U456 ( .B1(n619), .B2(n700), .A(n616), .ZN(n614) );
  NAND2_X4 U459 ( .A1(n700), .A2(n618), .ZN(n503) );
  NOR2_X4 U461 ( .A1(n1285), .A2(n1294), .ZN(n617) );
  NAND2_X4 U462 ( .A1(n1285), .A2(n1294), .ZN(n618) );
  XOR2_X2 U463 ( .A(n622), .B(n504), .Z(product[16]) );
  NAND2_X4 U465 ( .A1(n701), .A2(n621), .ZN(n504) );
  NOR2_X4 U467 ( .A1(n1295), .A2(n1304), .ZN(n620) );
  NAND2_X4 U468 ( .A1(n1295), .A2(n1304), .ZN(n621) );
  AOI21_X4 U470 ( .B1(n627), .B2(n702), .A(n624), .ZN(n622) );
  NAND2_X4 U473 ( .A1(n702), .A2(n626), .ZN(n505) );
  NOR2_X4 U475 ( .A1(n1305), .A2(n1314), .ZN(n625) );
  NAND2_X4 U476 ( .A1(n1305), .A2(n1314), .ZN(n626) );
  NAND2_X4 U479 ( .A1(n703), .A2(n629), .ZN(n506) );
  NOR2_X4 U481 ( .A1(n1315), .A2(n1322), .ZN(n628) );
  NAND2_X4 U482 ( .A1(n1315), .A2(n1322), .ZN(n629) );
  AOI21_X4 U484 ( .B1(n635), .B2(n704), .A(n632), .ZN(n630) );
  NAND2_X4 U487 ( .A1(n704), .A2(n634), .ZN(n507) );
  NOR2_X4 U489 ( .A1(n1323), .A2(n1330), .ZN(n633) );
  NAND2_X4 U490 ( .A1(n1323), .A2(n1330), .ZN(n634) );
  NAND2_X4 U493 ( .A1(n705), .A2(n637), .ZN(n508) );
  NOR2_X4 U495 ( .A1(n1331), .A2(n1338), .ZN(n636) );
  NAND2_X4 U496 ( .A1(n1331), .A2(n1338), .ZN(n637) );
  NAND2_X4 U501 ( .A1(n706), .A2(n642), .ZN(n509) );
  NOR2_X4 U503 ( .A1(n1339), .A2(n1344), .ZN(n641) );
  NAND2_X4 U504 ( .A1(n1339), .A2(n1344), .ZN(n642) );
  NAND2_X4 U507 ( .A1(n707), .A2(n645), .ZN(n510) );
  NOR2_X4 U509 ( .A1(n1345), .A2(n1350), .ZN(n644) );
  NAND2_X4 U510 ( .A1(n1345), .A2(n1350), .ZN(n645) );
  NAND2_X4 U515 ( .A1(n708), .A2(n650), .ZN(n511) );
  XOR2_X2 U519 ( .A(n654), .B(n512), .Z(product[8]) );
  NAND2_X4 U521 ( .A1(n709), .A2(n653), .ZN(n512) );
  NOR2_X4 U523 ( .A1(n1357), .A2(n1360), .ZN(n652) );
  NAND2_X4 U524 ( .A1(n1357), .A2(n1360), .ZN(n653) );
  AOI21_X4 U526 ( .B1(n710), .B2(n659), .A(n656), .ZN(n654) );
  NAND2_X4 U529 ( .A1(n710), .A2(n658), .ZN(n513) );
  NOR2_X4 U531 ( .A1(n1361), .A2(n1364), .ZN(n657) );
  NAND2_X4 U532 ( .A1(n1361), .A2(n1364), .ZN(n658) );
  XOR2_X2 U533 ( .A(n514), .B(n662), .Z(product[6]) );
  NAND2_X4 U535 ( .A1(n711), .A2(n661), .ZN(n514) );
  NOR2_X4 U537 ( .A1(n1365), .A2(n2087), .ZN(n660) );
  NAND2_X4 U538 ( .A1(n1365), .A2(n2087), .ZN(n661) );
  AOI21_X4 U540 ( .B1(n712), .B2(n667), .A(n664), .ZN(n662) );
  NAND2_X4 U543 ( .A1(n712), .A2(n666), .ZN(n515) );
  NOR2_X4 U545 ( .A1(n2088), .A2(n1369), .ZN(n665) );
  NAND2_X4 U546 ( .A1(n2088), .A2(n1369), .ZN(n666) );
  XOR2_X2 U547 ( .A(n516), .B(n670), .Z(product[4]) );
  NAND2_X4 U549 ( .A1(n713), .A2(n669), .ZN(n516) );
  NOR2_X4 U551 ( .A1(n1371), .A2(n2089), .ZN(n668) );
  NAND2_X4 U552 ( .A1(n1371), .A2(n2089), .ZN(n669) );
  XNOR2_X2 U553 ( .A(n517), .B(n675), .ZN(product[3]) );
  AOI21_X4 U554 ( .B1(n675), .B2(n714), .A(n672), .ZN(n670) );
  NAND2_X4 U557 ( .A1(n714), .A2(n674), .ZN(n517) );
  XOR2_X2 U561 ( .A(n676), .B(n677), .Z(product[2]) );
  NOR2_X4 U562 ( .A1(n676), .A2(n677), .ZN(n675) );
  XNOR2_X2 U564 ( .A(n679), .B(n680), .ZN(product[1]) );
  NAND2_X4 U565 ( .A1(n678), .A2(n680), .ZN(n677) );
  FA_X1 U576 ( .A(n1721), .B(n1745), .CI(n723), .CO(n719), .S(n720) );
  FA_X1 U577 ( .A(n727), .B(n1722), .CI(n1746), .CO(n721), .S(n722) );
  FA_X1 U579 ( .A(n1747), .B(n727), .CI(n730), .CO(n725), .S(n726) );
  FA_X1 U581 ( .A(n734), .B(n1748), .CI(n731), .CO(n728), .S(n729) );
  FA_X1 U582 ( .A(n736), .B(n1779), .CI(n1723), .CO(n730), .S(n731) );
  FA_X1 U583 ( .A(n740), .B(n1749), .CI(n735), .CO(n732), .S(n733) );
  FA_X1 U584 ( .A(n742), .B(n1724), .CI(n1780), .CO(n734), .S(n735) );
  FA_X1 U586 ( .A(n741), .B(n747), .CI(n745), .CO(n738), .S(n739) );
  FA_X1 U587 ( .A(n1781), .B(n742), .CI(n1750), .CO(n740), .S(n741) );
  FA_X1 U589 ( .A(n751), .B(n748), .CI(n746), .CO(n743), .S(n744) );
  FA_X1 U590 ( .A(n1751), .B(n1782), .CI(n753), .CO(n745), .S(n746) );
  FA_X1 U591 ( .A(n755), .B(n1814), .CI(n1725), .CO(n747), .S(n748) );
  FA_X1 U592 ( .A(n759), .B(n754), .CI(n752), .CO(n749), .S(n750) );
  FA_X1 U593 ( .A(n1752), .B(n1783), .CI(n761), .CO(n751), .S(n752) );
  FA_X1 U594 ( .A(n763), .B(n1726), .CI(n1815), .CO(n753), .S(n754) );
  FA_X1 U596 ( .A(n766), .B(n762), .CI(n760), .CO(n757), .S(n758) );
  FA_X1 U597 ( .A(n770), .B(n1753), .CI(n768), .CO(n759), .S(n760) );
  FA_X1 U598 ( .A(n1816), .B(n763), .CI(n1784), .CO(n761), .S(n762) );
  FA_X1 U600 ( .A(n774), .B(n769), .CI(n767), .CO(n764), .S(n765) );
  FA_X1 U601 ( .A(n771), .B(n778), .CI(n776), .CO(n766), .S(n767) );
  FA_X1 U602 ( .A(n1785), .B(n1754), .CI(n1817), .CO(n768), .S(n769) );
  FA_X1 U603 ( .A(n780), .B(n1849), .CI(n1727), .CO(n770), .S(n771) );
  FA_X1 U604 ( .A(n784), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U605 ( .A(n779), .B(n788), .CI(n786), .CO(n774), .S(n775) );
  FA_X1 U606 ( .A(n1786), .B(n1755), .CI(n1818), .CO(n776), .S(n777) );
  FA_X1 U607 ( .A(n790), .B(n1728), .CI(n1850), .CO(n778), .S(n779) );
  FA_X1 U609 ( .A(n793), .B(n787), .CI(n785), .CO(n782), .S(n783) );
  FA_X1 U610 ( .A(n789), .B(n797), .CI(n795), .CO(n784), .S(n785) );
  FA_X1 U611 ( .A(n1787), .B(n1819), .CI(n799), .CO(n786), .S(n787) );
  FA_X1 U612 ( .A(n1851), .B(n790), .CI(n1756), .CO(n788), .S(n789) );
  FA_X1 U614 ( .A(n803), .B(n796), .CI(n794), .CO(n791), .S(n792) );
  FA_X1 U615 ( .A(n798), .B(n807), .CI(n805), .CO(n793), .S(n794) );
  FA_X1 U616 ( .A(n809), .B(n1820), .CI(n800), .CO(n795), .S(n796) );
  FA_X1 U617 ( .A(n1852), .B(n1757), .CI(n1788), .CO(n797), .S(n798) );
  FA_X1 U618 ( .A(n811), .B(n1884), .CI(n1729), .CO(n799), .S(n800) );
  FA_X1 U619 ( .A(n815), .B(n806), .CI(n804), .CO(n801), .S(n802) );
  FA_X1 U620 ( .A(n808), .B(n819), .CI(n817), .CO(n803), .S(n804) );
  FA_X1 U621 ( .A(n821), .B(n1758), .CI(n810), .CO(n805), .S(n806) );
  FA_X1 U622 ( .A(n1853), .B(n1789), .CI(n1821), .CO(n807), .S(n808) );
  FA_X1 U623 ( .A(n823), .B(n1730), .CI(n1885), .CO(n809), .S(n810) );
  FA_X1 U625 ( .A(n826), .B(n818), .CI(n816), .CO(n813), .S(n814) );
  FA_X1 U626 ( .A(n820), .B(n822), .CI(n828), .CO(n815), .S(n816) );
  FA_X1 U627 ( .A(n832), .B(n1759), .CI(n830), .CO(n817), .S(n818) );
  FA_X1 U628 ( .A(n1822), .B(n1790), .CI(n1854), .CO(n819), .S(n820) );
  FA_X1 U629 ( .A(n834), .B(n823), .CI(n1886), .CO(n821), .S(n822) );
  FA_X1 U631 ( .A(n838), .B(n829), .CI(n827), .CO(n824), .S(n825) );
  FA_X1 U632 ( .A(n842), .B(n833), .CI(n840), .CO(n826), .S(n827) );
  FA_X1 U633 ( .A(n844), .B(n846), .CI(n831), .CO(n828), .S(n829) );
  FA_X1 U634 ( .A(n1823), .B(n1760), .CI(n1887), .CO(n830), .S(n831) );
  FA_X1 U635 ( .A(n1855), .B(n1791), .CI(n835), .CO(n832), .S(n833) );
  FA_X1 U636 ( .A(n848), .B(n1919), .CI(n1731), .CO(n834), .S(n835) );
  FA_X1 U637 ( .A(n852), .B(n841), .CI(n839), .CO(n836), .S(n837) );
  FA_X1 U638 ( .A(n843), .B(n856), .CI(n854), .CO(n838), .S(n839) );
  FA_X1 U639 ( .A(n858), .B(n847), .CI(n845), .CO(n840), .S(n841) );
  FA_X1 U640 ( .A(n1761), .B(n1824), .CI(n860), .CO(n842), .S(n843) );
  FA_X1 U641 ( .A(n1888), .B(n1792), .CI(n1856), .CO(n844), .S(n845) );
  FA_X1 U642 ( .A(n1732), .B(n862), .CI(n1920), .CO(n846), .S(n847) );
  FA_X1 U644 ( .A(n865), .B(n855), .CI(n853), .CO(n850), .S(n851) );
  FA_X1 U645 ( .A(n857), .B(n869), .CI(n867), .CO(n852), .S(n853) );
  FA_X1 U646 ( .A(n861), .B(n871), .CI(n859), .CO(n854), .S(n855) );
  FA_X1 U647 ( .A(n1857), .B(n1762), .CI(n873), .CO(n856), .S(n857) );
  FA_X1 U648 ( .A(n1889), .B(n1793), .CI(n875), .CO(n858), .S(n859) );
  FA_X1 U649 ( .A(n1921), .B(n862), .CI(n1825), .CO(n860), .S(n861) );
  FA_X1 U651 ( .A(n879), .B(n868), .CI(n866), .CO(n863), .S(n864) );
  FA_X1 U652 ( .A(n870), .B(n883), .CI(n881), .CO(n865), .S(n866) );
  FA_X1 U653 ( .A(n874), .B(n885), .CI(n872), .CO(n867), .S(n868) );
  FA_X1 U654 ( .A(n889), .B(n876), .CI(n887), .CO(n869), .S(n870) );
  FA_X1 U655 ( .A(n1858), .B(n1922), .CI(n1890), .CO(n871), .S(n872) );
  FA_X1 U656 ( .A(n1826), .B(n1763), .CI(n1794), .CO(n873), .S(n874) );
  FA_X1 U657 ( .A(n891), .B(n3220), .CI(n1733), .CO(n875), .S(n876) );
  FA_X1 U658 ( .A(n895), .B(n882), .CI(n880), .CO(n877), .S(n878) );
  FA_X1 U659 ( .A(n884), .B(n899), .CI(n897), .CO(n879), .S(n880) );
  FA_X1 U660 ( .A(n888), .B(n901), .CI(n886), .CO(n881), .S(n882) );
  FA_X1 U661 ( .A(n890), .B(n905), .CI(n903), .CO(n883), .S(n884) );
  FA_X1 U662 ( .A(n1891), .B(n1859), .CI(n1923), .CO(n885), .S(n886) );
  FA_X1 U663 ( .A(n1827), .B(n1764), .CI(n1795), .CO(n887), .S(n888) );
  FA_X1 U664 ( .A(n907), .B(n892), .CI(n1955), .CO(n889), .S(n890) );
  FA_X1 U666 ( .A(n911), .B(n898), .CI(n896), .CO(n893), .S(n894) );
  FA_X1 U667 ( .A(n900), .B(n915), .CI(n913), .CO(n895), .S(n896) );
  FA_X1 U668 ( .A(n904), .B(n917), .CI(n902), .CO(n897), .S(n898) );
  FA_X1 U669 ( .A(n921), .B(n906), .CI(n919), .CO(n899), .S(n900) );
  FA_X1 U670 ( .A(n1892), .B(n1796), .CI(n1924), .CO(n901), .S(n902) );
  FA_X1 U671 ( .A(n1828), .B(n1956), .CI(n1860), .CO(n903), .S(n904) );
  FA_X1 U672 ( .A(n908), .B(n1734), .CI(n923), .CO(n905), .S(n906) );
  FA_X1 U674 ( .A(n927), .B(n914), .CI(n912), .CO(n909), .S(n910) );
  FA_X1 U675 ( .A(n916), .B(n931), .CI(n929), .CO(n911), .S(n912) );
  FA_X1 U676 ( .A(n920), .B(n933), .CI(n918), .CO(n913), .S(n914) );
  FA_X1 U677 ( .A(n935), .B(n937), .CI(n922), .CO(n915), .S(n916) );
  FA_X1 U678 ( .A(n1893), .B(n1829), .CI(n1957), .CO(n917), .S(n918) );
  FA_X1 U679 ( .A(n1925), .B(n1861), .CI(n939), .CO(n919), .S(n920) );
  FA_X1 U680 ( .A(n1765), .B(n1797), .CI(n924), .CO(n921), .S(n922) );
  FA_X1 U681 ( .A(n941), .B(n1989), .CI(n1735), .CO(n923), .S(n924) );
  FA_X1 U682 ( .A(n945), .B(n930), .CI(n928), .CO(n925), .S(n926) );
  FA_X1 U683 ( .A(n932), .B(n949), .CI(n947), .CO(n927), .S(n928) );
  FA_X1 U684 ( .A(n951), .B(n936), .CI(n934), .CO(n929), .S(n930) );
  FA_X1 U685 ( .A(n953), .B(n955), .CI(n938), .CO(n931), .S(n932) );
  FA_X1 U686 ( .A(n957), .B(n1894), .CI(n940), .CO(n933), .S(n934) );
  FA_X1 U687 ( .A(n1926), .B(n1830), .CI(n1958), .CO(n935), .S(n936) );
  FA_X1 U688 ( .A(n1798), .B(n1990), .CI(n1862), .CO(n937), .S(n938) );
  FA_X1 U689 ( .A(n1736), .B(n959), .CI(n1766), .CO(n939), .S(n940) );
  FA_X1 U691 ( .A(n962), .B(n948), .CI(n946), .CO(n943), .S(n944) );
  FA_X1 U692 ( .A(n950), .B(n966), .CI(n964), .CO(n945), .S(n946) );
  FA_X1 U693 ( .A(n968), .B(n954), .CI(n952), .CO(n947), .S(n948) );
  FA_X1 U694 ( .A(n970), .B(n972), .CI(n956), .CO(n949), .S(n950) );
  FA_X1 U695 ( .A(n974), .B(n1895), .CI(n958), .CO(n951), .S(n952) );
  FA_X1 U696 ( .A(n1927), .B(n1831), .CI(n1959), .CO(n953), .S(n954) );
  FA_X1 U697 ( .A(n1767), .B(n1991), .CI(n1863), .CO(n955), .S(n956) );
  FA_X1 U698 ( .A(n1799), .B(n959), .CI(n976), .CO(n957), .S(n958) );
  FA_X1 U700 ( .A(n980), .B(n965), .CI(n963), .CO(n960), .S(n961) );
  FA_X1 U701 ( .A(n967), .B(n969), .CI(n982), .CO(n962), .S(n963) );
  FA_X1 U702 ( .A(n986), .B(n971), .CI(n984), .CO(n964), .S(n965) );
  FA_X1 U703 ( .A(n975), .B(n988), .CI(n973), .CO(n966), .S(n967) );
  FA_X1 U704 ( .A(n992), .B(n1960), .CI(n990), .CO(n968), .S(n969) );
  FA_X1 U705 ( .A(n1928), .B(n1992), .CI(n994), .CO(n970), .S(n971) );
  FA_X1 U706 ( .A(n1896), .B(n977), .CI(n1864), .CO(n972), .S(n973) );
  FA_X1 U707 ( .A(n1832), .B(n1768), .CI(n1800), .CO(n974), .S(n975) );
  FA_X1 U708 ( .A(n2024), .B(n2059), .CI(n1737), .CO(n976), .S(n977) );
  FA_X1 U709 ( .A(n998), .B(n983), .CI(n981), .CO(n978), .S(n979) );
  FA_X1 U710 ( .A(n985), .B(n987), .CI(n1000), .CO(n980), .S(n981) );
  FA_X1 U711 ( .A(n1004), .B(n989), .CI(n1002), .CO(n982), .S(n983) );
  FA_X1 U712 ( .A(n993), .B(n1006), .CI(n991), .CO(n984), .S(n985) );
  FA_X1 U713 ( .A(n1010), .B(n995), .CI(n1008), .CO(n986), .S(n987) );
  FA_X1 U714 ( .A(n1865), .B(n1929), .CI(n1961), .CO(n988), .S(n989) );
  FA_X1 U715 ( .A(n1897), .B(n1012), .CI(n1993), .CO(n990), .S(n991) );
  FA_X1 U716 ( .A(n2025), .B(n1769), .CI(n1833), .CO(n992), .S(n993) );
  FA_X1 U717 ( .A(n1738), .B(n262), .CI(n1801), .CO(n994), .S(n995) );
  FA_X1 U718 ( .A(n1016), .B(n1001), .CI(n999), .CO(n996), .S(n997) );
  FA_X1 U719 ( .A(n1003), .B(n1005), .CI(n1018), .CO(n998), .S(n999) );
  FA_X1 U720 ( .A(n1022), .B(n1009), .CI(n1020), .CO(n1000), .S(n1001) );
  FA_X1 U721 ( .A(n1011), .B(n1024), .CI(n1007), .CO(n1002), .S(n1003) );
  FA_X1 U722 ( .A(n1028), .B(n1013), .CI(n1026), .CO(n1004), .S(n1005) );
  FA_X1 U723 ( .A(n1866), .B(n1930), .CI(n1962), .CO(n1006), .S(n1007) );
  FA_X1 U724 ( .A(n1994), .B(n1898), .CI(n1030), .CO(n1008), .S(n1009) );
  FA_X1 U725 ( .A(n2026), .B(n1834), .CI(n1802), .CO(n1010), .S(n1011) );
  FA_X1 U726 ( .A(n1739), .B(n262), .CI(n1770), .CO(n1012), .S(n1013) );
  FA_X1 U727 ( .A(n1034), .B(n1019), .CI(n1017), .CO(n1014), .S(n1015) );
  FA_X1 U728 ( .A(n1021), .B(n1023), .CI(n1036), .CO(n1016), .S(n1017) );
  FA_X1 U729 ( .A(n1040), .B(n1027), .CI(n1038), .CO(n1018), .S(n1019) );
  FA_X1 U730 ( .A(n1029), .B(n1042), .CI(n1025), .CO(n1020), .S(n1021) );
  FA_X1 U731 ( .A(n1046), .B(n1031), .CI(n1044), .CO(n1022), .S(n1023) );
  FA_X1 U732 ( .A(n1963), .B(n1899), .CI(n1995), .CO(n1024), .S(n1025) );
  FA_X1 U733 ( .A(n2027), .B(n1931), .CI(n1048), .CO(n1026), .S(n1027) );
  FA_X1 U734 ( .A(n1867), .B(n1803), .CI(n1835), .CO(n1028), .S(n1029) );
  FA_X1 U735 ( .A(n1740), .B(n262), .CI(n1771), .CO(n1030), .S(n1031) );
  FA_X1 U736 ( .A(n1052), .B(n1037), .CI(n1035), .CO(n1032), .S(n1033) );
  FA_X1 U737 ( .A(n1039), .B(n1041), .CI(n1054), .CO(n1034), .S(n1035) );
  FA_X1 U738 ( .A(n1058), .B(n1045), .CI(n1056), .CO(n1036), .S(n1037) );
  FA_X1 U739 ( .A(n1047), .B(n1060), .CI(n1043), .CO(n1038), .S(n1039) );
  FA_X1 U740 ( .A(n1064), .B(n1049), .CI(n1062), .CO(n1040), .S(n1041) );
  FA_X1 U741 ( .A(n1900), .B(n1964), .CI(n1066), .CO(n1042), .S(n1043) );
  FA_X1 U742 ( .A(n2028), .B(n1932), .CI(n1996), .CO(n1044), .S(n1045) );
  FA_X1 U743 ( .A(n2060), .B(n1836), .CI(n1868), .CO(n1046), .S(n1047) );
  FA_X1 U744 ( .A(n1772), .B(n1741), .CI(n1804), .CO(n1048), .S(n1049) );
  FA_X1 U745 ( .A(n1070), .B(n1055), .CI(n1053), .CO(n1050), .S(n1051) );
  FA_X1 U746 ( .A(n1057), .B(n1059), .CI(n1072), .CO(n1052), .S(n1053) );
  FA_X1 U747 ( .A(n1076), .B(n1063), .CI(n1074), .CO(n1054), .S(n1055) );
  FA_X1 U748 ( .A(n1065), .B(n1078), .CI(n1061), .CO(n1056), .S(n1057) );
  FA_X1 U749 ( .A(n1067), .B(n1082), .CI(n1080), .CO(n1058), .S(n1059) );
  FA_X1 U750 ( .A(n1933), .B(n1965), .CI(n1997), .CO(n1060), .S(n1061) );
  FA_X1 U751 ( .A(n2029), .B(n1901), .CI(n1084), .CO(n1062), .S(n1063) );
  FA_X1 U752 ( .A(n2061), .B(n1869), .CI(n1837), .CO(n1064), .S(n1065) );
  FA_X1 U753 ( .A(n1773), .B(n1742), .CI(n1805), .CO(n1066), .S(n1067) );
  FA_X1 U754 ( .A(n1088), .B(n1073), .CI(n1071), .CO(n1068), .S(n1069) );
  FA_X1 U755 ( .A(n1075), .B(n1092), .CI(n1090), .CO(n1070), .S(n1071) );
  FA_X1 U756 ( .A(n1079), .B(n1094), .CI(n1077), .CO(n1072), .S(n1073) );
  FA_X1 U757 ( .A(n1096), .B(n1098), .CI(n1081), .CO(n1074), .S(n1075) );
  FA_X1 U758 ( .A(n1085), .B(n1100), .CI(n1083), .CO(n1076), .S(n1077) );
  FA_X1 U759 ( .A(n1998), .B(n2062), .CI(n2030), .CO(n1078), .S(n1079) );
  FA_X1 U760 ( .A(n1966), .B(n1870), .CI(n1934), .CO(n1080), .S(n1081) );
  FA_X1 U761 ( .A(n1102), .B(n1838), .CI(n1902), .CO(n1082), .S(n1083) );
  FA_X1 U762 ( .A(n1774), .B(n1743), .CI(n1806), .CO(n1084), .S(n1085) );
  FA_X1 U763 ( .A(n1106), .B(n1091), .CI(n1089), .CO(n1086), .S(n1087) );
  FA_X1 U764 ( .A(n1108), .B(n1110), .CI(n1093), .CO(n1088), .S(n1089) );
  FA_X1 U765 ( .A(n1097), .B(n1099), .CI(n1095), .CO(n1090), .S(n1091) );
  FA_X1 U766 ( .A(n1114), .B(n1116), .CI(n1112), .CO(n1092), .S(n1093) );
  FA_X1 U767 ( .A(n1118), .B(n1999), .CI(n1101), .CO(n1094), .S(n1095) );
  FA_X1 U768 ( .A(n2063), .B(n1935), .CI(n2031), .CO(n1096), .S(n1097) );
  FA_X1 U769 ( .A(n1903), .B(n1103), .CI(n1967), .CO(n1098), .S(n1099) );
  FA_X1 U770 ( .A(n1871), .B(n1807), .CI(n1839), .CO(n1100), .S(n1101) );
  FA_X1 U771 ( .A(n1775), .B(n1744), .CI(n1120), .CO(n1102), .S(n1103) );
  FA_X1 U772 ( .A(n1124), .B(n1109), .CI(n1107), .CO(n1104), .S(n1105) );
  FA_X1 U773 ( .A(n1126), .B(n1128), .CI(n1111), .CO(n1106), .S(n1107) );
  FA_X1 U774 ( .A(n1115), .B(n1117), .CI(n1113), .CO(n1108), .S(n1109) );
  FA_X1 U775 ( .A(n1132), .B(n1119), .CI(n1130), .CO(n1110), .S(n1111) );
  FA_X1 U776 ( .A(n2064), .B(n2000), .CI(n1134), .CO(n1112), .S(n1113) );
  FA_X1 U777 ( .A(n2032), .B(n1936), .CI(n1136), .CO(n1114), .S(n1115) );
  FA_X1 U778 ( .A(n1872), .B(n1904), .CI(n1968), .CO(n1116), .S(n1117) );
  FA_X1 U779 ( .A(n1808), .B(n1121), .CI(n1840), .CO(n1118), .S(n1119) );
  HA_X1 U780 ( .A(n1776), .B(n1138), .CO(n1120), .S(n1121) );
  FA_X1 U781 ( .A(n1142), .B(n1127), .CI(n1125), .CO(n1122), .S(n1123) );
  FA_X1 U782 ( .A(n1129), .B(n1146), .CI(n1144), .CO(n1124), .S(n1125) );
  FA_X1 U783 ( .A(n1133), .B(n1148), .CI(n1131), .CO(n1126), .S(n1127) );
  FA_X1 U784 ( .A(n1135), .B(n1137), .CI(n1150), .CO(n1128), .S(n1129) );
  FA_X1 U785 ( .A(n2033), .B(n2065), .CI(n1152), .CO(n1130), .S(n1131) );
  FA_X1 U786 ( .A(n2001), .B(n1905), .CI(n1969), .CO(n1132), .S(n1133) );
  FA_X1 U787 ( .A(n1154), .B(n1873), .CI(n1937), .CO(n1134), .S(n1135) );
  FA_X1 U788 ( .A(n1139), .B(n1809), .CI(n1841), .CO(n1136), .S(n1137) );
  HA_X1 U789 ( .A(n1156), .B(n1777), .CO(n1138), .S(n1139) );
  FA_X1 U790 ( .A(n1160), .B(n1145), .CI(n1143), .CO(n1140), .S(n1141) );
  FA_X1 U791 ( .A(n1147), .B(n1149), .CI(n1162), .CO(n1142), .S(n1143) );
  FA_X1 U792 ( .A(n1164), .B(n1166), .CI(n1151), .CO(n1144), .S(n1145) );
  FA_X1 U793 ( .A(n1153), .B(n2002), .CI(n1168), .CO(n1146), .S(n1147) );
  FA_X1 U794 ( .A(n1170), .B(n2034), .CI(n2066), .CO(n1148), .S(n1149) );
  FA_X1 U795 ( .A(n1938), .B(n1155), .CI(n1970), .CO(n1150), .S(n1151) );
  FA_X1 U796 ( .A(n1874), .B(n1842), .CI(n1906), .CO(n1152), .S(n1153) );
  FA_X1 U797 ( .A(n1810), .B(n1157), .CI(n1172), .CO(n1154), .S(n1155) );
  HA_X1 U798 ( .A(n289), .B(n1778), .CO(n1156), .S(n1157) );
  FA_X1 U799 ( .A(n1176), .B(n1163), .CI(n1161), .CO(n1158), .S(n1159) );
  FA_X1 U800 ( .A(n1165), .B(n1167), .CI(n1178), .CO(n1160), .S(n1161) );
  FA_X1 U801 ( .A(n1169), .B(n1182), .CI(n1180), .CO(n1162), .S(n1163) );
  FA_X1 U802 ( .A(n1184), .B(n2003), .CI(n1171), .CO(n1164), .S(n1165) );
  FA_X1 U803 ( .A(n2067), .B(n2035), .CI(n1186), .CO(n1166), .S(n1167) );
  FA_X1 U804 ( .A(n1907), .B(n1939), .CI(n1971), .CO(n1168), .S(n1169) );
  FA_X1 U805 ( .A(n1843), .B(n1173), .CI(n1875), .CO(n1170), .S(n1171) );
  HA_X1 U806 ( .A(n1811), .B(n1188), .CO(n1172), .S(n1173) );
  FA_X1 U807 ( .A(n1192), .B(n1179), .CI(n1177), .CO(n1174), .S(n1175) );
  FA_X1 U808 ( .A(n1181), .B(n1183), .CI(n1194), .CO(n1176), .S(n1177) );
  FA_X1 U809 ( .A(n1198), .B(n1185), .CI(n1196), .CO(n1178), .S(n1179) );
  FA_X1 U810 ( .A(n1200), .B(n2068), .CI(n1187), .CO(n1180), .S(n1181) );
  FA_X1 U811 ( .A(n2004), .B(n1940), .CI(n2036), .CO(n1182), .S(n1183) );
  FA_X1 U812 ( .A(n1202), .B(n1908), .CI(n1972), .CO(n1184), .S(n1185) );
  FA_X1 U813 ( .A(n1189), .B(n1844), .CI(n1876), .CO(n1186), .S(n1187) );
  HA_X1 U814 ( .A(n1204), .B(n1812), .CO(n1188), .S(n1189) );
  FA_X1 U815 ( .A(n1208), .B(n1195), .CI(n1193), .CO(n1190), .S(n1191) );
  FA_X1 U816 ( .A(n1197), .B(n1199), .CI(n1210), .CO(n1192), .S(n1193) );
  FA_X1 U817 ( .A(n1214), .B(n1201), .CI(n1212), .CO(n1194), .S(n1195) );
  FA_X1 U818 ( .A(n2037), .B(n2069), .CI(n1216), .CO(n1196), .S(n1197) );
  FA_X1 U819 ( .A(n1973), .B(n1203), .CI(n2005), .CO(n1198), .S(n1199) );
  FA_X1 U820 ( .A(n1941), .B(n1877), .CI(n1909), .CO(n1200), .S(n1201) );
  FA_X1 U821 ( .A(n1845), .B(n1205), .CI(n1218), .CO(n1202), .S(n1203) );
  HA_X1 U822 ( .A(n286), .B(n1813), .CO(n1204), .S(n1205) );
  FA_X1 U823 ( .A(n1222), .B(n1211), .CI(n1209), .CO(n1206), .S(n1207) );
  FA_X1 U824 ( .A(n1213), .B(n1215), .CI(n1224), .CO(n1208), .S(n1209) );
  FA_X1 U825 ( .A(n1217), .B(n1228), .CI(n1226), .CO(n1210), .S(n1211) );
  FA_X1 U826 ( .A(n2038), .B(n2070), .CI(n1230), .CO(n1212), .S(n1213) );
  FA_X1 U827 ( .A(n1942), .B(n1974), .CI(n2006), .CO(n1214), .S(n1215) );
  FA_X1 U828 ( .A(n1878), .B(n1219), .CI(n1910), .CO(n1216), .S(n1217) );
  HA_X1 U829 ( .A(n1846), .B(n1232), .CO(n1218), .S(n1219) );
  FA_X1 U830 ( .A(n1236), .B(n1225), .CI(n1223), .CO(n1220), .S(n1221) );
  FA_X1 U831 ( .A(n1227), .B(n1240), .CI(n1238), .CO(n1222), .S(n1223) );
  FA_X1 U832 ( .A(n1231), .B(n1242), .CI(n1229), .CO(n1224), .S(n1225) );
  FA_X1 U833 ( .A(n2071), .B(n1975), .CI(n2039), .CO(n1226), .S(n1227) );
  FA_X1 U834 ( .A(n1244), .B(n1943), .CI(n2007), .CO(n1228), .S(n1229) );
  FA_X1 U835 ( .A(n1233), .B(n1879), .CI(n1911), .CO(n1230), .S(n1231) );
  HA_X1 U836 ( .A(n1246), .B(n1847), .CO(n1232), .S(n1233) );
  FA_X1 U837 ( .A(n1250), .B(n1239), .CI(n1237), .CO(n1234), .S(n1235) );
  FA_X1 U838 ( .A(n1252), .B(n1254), .CI(n1241), .CO(n1236), .S(n1237) );
  FA_X1 U839 ( .A(n1256), .B(n2040), .CI(n1243), .CO(n1238), .S(n1239) );
  FA_X1 U840 ( .A(n2008), .B(n1245), .CI(n2072), .CO(n1240), .S(n1241) );
  FA_X1 U841 ( .A(n1944), .B(n1912), .CI(n1976), .CO(n1242), .S(n1243) );
  FA_X1 U842 ( .A(n1880), .B(n1247), .CI(n1258), .CO(n1244), .S(n1245) );
  HA_X1 U843 ( .A(n283), .B(n1848), .CO(n1246), .S(n1247) );
  FA_X1 U844 ( .A(n1262), .B(n1253), .CI(n1251), .CO(n1248), .S(n1249) );
  FA_X1 U845 ( .A(n1264), .B(n1257), .CI(n1255), .CO(n1250), .S(n1251) );
  FA_X1 U846 ( .A(n1268), .B(n2041), .CI(n1266), .CO(n1252), .S(n1253) );
  FA_X1 U847 ( .A(n1977), .B(n2009), .CI(n2073), .CO(n1254), .S(n1255) );
  FA_X1 U848 ( .A(n1913), .B(n1259), .CI(n1945), .CO(n1256), .S(n1257) );
  HA_X1 U849 ( .A(n1881), .B(n1270), .CO(n1258), .S(n1259) );
  FA_X1 U850 ( .A(n1274), .B(n1265), .CI(n1263), .CO(n1260), .S(n1261) );
  FA_X1 U851 ( .A(n1267), .B(n1269), .CI(n1276), .CO(n1262), .S(n1263) );
  FA_X1 U852 ( .A(n2074), .B(n2010), .CI(n1278), .CO(n1264), .S(n1265) );
  FA_X1 U853 ( .A(n1280), .B(n1978), .CI(n2042), .CO(n1266), .S(n1267) );
  FA_X1 U854 ( .A(n1271), .B(n1914), .CI(n1946), .CO(n1268), .S(n1269) );
  HA_X1 U855 ( .A(n1282), .B(n1882), .CO(n1270), .S(n1271) );
  FA_X1 U856 ( .A(n1277), .B(n1286), .CI(n1275), .CO(n1272), .S(n1273) );
  FA_X1 U857 ( .A(n1279), .B(n1290), .CI(n1288), .CO(n1274), .S(n1275) );
  FA_X1 U858 ( .A(n2043), .B(n1281), .CI(n2075), .CO(n1276), .S(n1277) );
  FA_X1 U859 ( .A(n2011), .B(n1947), .CI(n1979), .CO(n1278), .S(n1279) );
  FA_X1 U860 ( .A(n1915), .B(n1283), .CI(n1292), .CO(n1280), .S(n1281) );
  HA_X1 U861 ( .A(n280), .B(n1883), .CO(n1282), .S(n1283) );
  FA_X1 U862 ( .A(n1296), .B(n1289), .CI(n1287), .CO(n1284), .S(n1285) );
  FA_X1 U863 ( .A(n1298), .B(n1300), .CI(n1291), .CO(n1286), .S(n1287) );
  FA_X1 U864 ( .A(n2012), .B(n2044), .CI(n2076), .CO(n1288), .S(n1289) );
  FA_X1 U865 ( .A(n1948), .B(n1293), .CI(n1980), .CO(n1290), .S(n1291) );
  HA_X1 U866 ( .A(n1916), .B(n1302), .CO(n1292), .S(n1293) );
  FA_X1 U867 ( .A(n1306), .B(n1299), .CI(n1297), .CO(n1294), .S(n1295) );
  FA_X1 U868 ( .A(n1308), .B(n2045), .CI(n1301), .CO(n1296), .S(n1297) );
  FA_X1 U869 ( .A(n1310), .B(n2013), .CI(n2077), .CO(n1298), .S(n1299) );
  FA_X1 U870 ( .A(n1303), .B(n1949), .CI(n1981), .CO(n1300), .S(n1301) );
  HA_X1 U871 ( .A(n1312), .B(n1917), .CO(n1302), .S(n1303) );
  FA_X1 U872 ( .A(n1316), .B(n1309), .CI(n1307), .CO(n1304), .S(n1305) );
  FA_X1 U873 ( .A(n2078), .B(n1311), .CI(n1318), .CO(n1306), .S(n1307) );
  FA_X1 U874 ( .A(n2046), .B(n1982), .CI(n2014), .CO(n1308), .S(n1309) );
  FA_X1 U875 ( .A(n1950), .B(n1313), .CI(n1320), .CO(n1310), .S(n1311) );
  HA_X1 U876 ( .A(n277), .B(n1918), .CO(n1312), .S(n1313) );
  FA_X1 U877 ( .A(n1324), .B(n1319), .CI(n1317), .CO(n1314), .S(n1315) );
  FA_X1 U878 ( .A(n2047), .B(n2079), .CI(n1326), .CO(n1316), .S(n1317) );
  FA_X1 U879 ( .A(n1983), .B(n1321), .CI(n2015), .CO(n1318), .S(n1319) );
  HA_X1 U880 ( .A(n1951), .B(n1328), .CO(n1320), .S(n1321) );
  FA_X1 U881 ( .A(n1327), .B(n1332), .CI(n1325), .CO(n1322), .S(n1323) );
  FA_X1 U882 ( .A(n1334), .B(n2048), .CI(n2080), .CO(n1324), .S(n1325) );
  FA_X1 U883 ( .A(n1329), .B(n1984), .CI(n2016), .CO(n1326), .S(n1327) );
  HA_X1 U884 ( .A(n1336), .B(n1952), .CO(n1328), .S(n1329) );
  FA_X1 U885 ( .A(n1340), .B(n1335), .CI(n1333), .CO(n1330), .S(n1331) );
  FA_X1 U886 ( .A(n2081), .B(n2017), .CI(n2049), .CO(n1332), .S(n1333) );
  FA_X1 U887 ( .A(n1985), .B(n1337), .CI(n1342), .CO(n1334), .S(n1335) );
  HA_X1 U888 ( .A(n274), .B(n1953), .CO(n1336), .S(n1337) );
  FA_X1 U889 ( .A(n1346), .B(n2082), .CI(n1341), .CO(n1338), .S(n1339) );
  FA_X1 U890 ( .A(n2018), .B(n1343), .CI(n2050), .CO(n1340), .S(n1341) );
  HA_X1 U891 ( .A(n1986), .B(n1348), .CO(n1342), .S(n1343) );
  FA_X1 U892 ( .A(n1352), .B(n2083), .CI(n1347), .CO(n1344), .S(n1345) );
  FA_X1 U893 ( .A(n1349), .B(n2019), .CI(n2051), .CO(n1346), .S(n1347) );
  HA_X1 U894 ( .A(n1354), .B(n1987), .CO(n1348), .S(n1349) );
  FA_X1 U895 ( .A(n2084), .B(n2052), .CI(n1353), .CO(n1350), .S(n1351) );
  FA_X1 U896 ( .A(n2020), .B(n1355), .CI(n1358), .CO(n1352), .S(n1353) );
  HA_X1 U897 ( .A(n271), .B(n1988), .CO(n1354), .S(n1355) );
  FA_X1 U898 ( .A(n2053), .B(n1359), .CI(n2085), .CO(n1356), .S(n1357) );
  HA_X1 U899 ( .A(n2021), .B(n1362), .CO(n1358), .S(n1359) );
  FA_X1 U900 ( .A(n1363), .B(n2054), .CI(n2086), .CO(n1360), .S(n1361) );
  HA_X1 U901 ( .A(n1366), .B(n2022), .CO(n1362), .S(n1363) );
  FA_X1 U902 ( .A(n2055), .B(n1367), .CI(n1368), .CO(n1364), .S(n1365) );
  HA_X1 U903 ( .A(n268), .B(n2023), .CO(n1366), .S(n1367) );
  HA_X1 U904 ( .A(n2056), .B(n1370), .CO(n1368), .S(n1369) );
  HA_X1 U905 ( .A(n1372), .B(n2057), .CO(n1370), .S(n1371) );
  HA_X1 U906 ( .A(n265), .B(n2058), .CO(n1372), .S(n1373) );
  OAI21_X4 U907 ( .B1(n2808), .B2(n3157), .A(n2094), .ZN(n1720) );
  NAND2_X4 U908 ( .A1(n388), .A2(n484), .ZN(n2094) );
  OAI21_X4 U909 ( .B1(n2809), .B2(n3157), .A(n2095), .ZN(n717) );
  AOI21_X4 U910 ( .B1(n388), .B2(n481), .A(n1374), .ZN(n2095) );
  AND2_X4 U911 ( .A1(n333), .A2(n484), .ZN(n1374) );
  OAI21_X4 U912 ( .B1(n2810), .B2(n3157), .A(n2096), .ZN(n1721) );
  AOI222_X2 U913 ( .A1(n3145), .A2(n484), .B1(n333), .B2(n481), .C1(n388), 
        .C2(n478), .ZN(n2096) );
  OAI21_X4 U914 ( .B1(n2811), .B2(n3157), .A(n2097), .ZN(n1722) );
  AOI222_X2 U915 ( .A1(n3144), .A2(n481), .B1(n333), .B2(n478), .C1(n388), 
        .C2(n475), .ZN(n2097) );
  OAI21_X4 U916 ( .B1(n2812), .B2(n3157), .A(n2098), .ZN(n723) );
  AOI222_X2 U917 ( .A1(n3145), .A2(n478), .B1(n333), .B2(n475), .C1(n388), 
        .C2(n472), .ZN(n2098) );
  OAI21_X4 U918 ( .B1(n2813), .B2(n3157), .A(n2099), .ZN(n1723) );
  AOI222_X2 U919 ( .A1(n3144), .A2(n475), .B1(n333), .B2(n472), .C1(n388), 
        .C2(n469), .ZN(n2099) );
  OAI21_X4 U920 ( .B1(n2814), .B2(n3157), .A(n2100), .ZN(n1724) );
  AOI222_X2 U921 ( .A1(n3145), .A2(n472), .B1(n333), .B2(n469), .C1(n388), 
        .C2(n466), .ZN(n2100) );
  OAI21_X4 U922 ( .B1(n2815), .B2(n3157), .A(n2101), .ZN(n736) );
  AOI222_X2 U923 ( .A1(n3144), .A2(n469), .B1(n333), .B2(n466), .C1(n388), 
        .C2(n463), .ZN(n2101) );
  OAI21_X4 U924 ( .B1(n2816), .B2(n3157), .A(n2102), .ZN(n1725) );
  AOI222_X2 U925 ( .A1(n3145), .A2(n466), .B1(n333), .B2(n463), .C1(n388), 
        .C2(n460), .ZN(n2102) );
  OAI21_X4 U926 ( .B1(n2817), .B2(n3157), .A(n2103), .ZN(n1726) );
  AOI222_X2 U927 ( .A1(n3144), .A2(n463), .B1(n333), .B2(n460), .C1(n388), 
        .C2(n457), .ZN(n2103) );
  OAI21_X4 U928 ( .B1(n2818), .B2(n3157), .A(n2104), .ZN(n755) );
  AOI222_X2 U929 ( .A1(n3145), .A2(n460), .B1(n333), .B2(n457), .C1(n388), 
        .C2(n454), .ZN(n2104) );
  OAI21_X4 U930 ( .B1(n2819), .B2(n3157), .A(n2105), .ZN(n1727) );
  AOI222_X2 U931 ( .A1(n3144), .A2(n457), .B1(n333), .B2(n454), .C1(n388), 
        .C2(n451), .ZN(n2105) );
  OAI21_X4 U932 ( .B1(n2820), .B2(n3157), .A(n2106), .ZN(n1728) );
  AOI222_X2 U933 ( .A1(n3145), .A2(n454), .B1(n333), .B2(n451), .C1(n388), 
        .C2(n448), .ZN(n2106) );
  OAI21_X4 U934 ( .B1(n2821), .B2(n3157), .A(n2107), .ZN(n780) );
  AOI222_X2 U935 ( .A1(n3144), .A2(n451), .B1(n333), .B2(n448), .C1(n388), 
        .C2(n445), .ZN(n2107) );
  OAI21_X4 U936 ( .B1(n2822), .B2(n3157), .A(n2108), .ZN(n1729) );
  AOI222_X2 U937 ( .A1(n3145), .A2(n448), .B1(n333), .B2(n445), .C1(n388), 
        .C2(n442), .ZN(n2108) );
  OAI21_X4 U938 ( .B1(n2823), .B2(n3157), .A(n2109), .ZN(n1730) );
  AOI222_X2 U939 ( .A1(n3144), .A2(n445), .B1(n333), .B2(n442), .C1(n388), 
        .C2(n439), .ZN(n2109) );
  OAI21_X4 U940 ( .B1(n2824), .B2(n3157), .A(n2110), .ZN(n811) );
  AOI222_X2 U941 ( .A1(n3145), .A2(n442), .B1(n333), .B2(n439), .C1(n388), 
        .C2(n436), .ZN(n2110) );
  OAI21_X4 U942 ( .B1(n2825), .B2(n3157), .A(n2111), .ZN(n1731) );
  AOI222_X2 U943 ( .A1(n3144), .A2(n439), .B1(n333), .B2(n436), .C1(n388), 
        .C2(n433), .ZN(n2111) );
  OAI21_X4 U944 ( .B1(n2826), .B2(n3157), .A(n2112), .ZN(n1732) );
  AOI222_X2 U945 ( .A1(n3145), .A2(n436), .B1(n333), .B2(n433), .C1(n388), 
        .C2(n430), .ZN(n2112) );
  OAI21_X4 U946 ( .B1(n2827), .B2(n3157), .A(n2113), .ZN(n848) );
  AOI222_X2 U947 ( .A1(n3144), .A2(n433), .B1(n333), .B2(n430), .C1(n388), 
        .C2(n427), .ZN(n2113) );
  OAI21_X4 U948 ( .B1(n2828), .B2(n3157), .A(n2114), .ZN(n1733) );
  AOI222_X2 U949 ( .A1(n3145), .A2(n430), .B1(n333), .B2(n427), .C1(n388), 
        .C2(n424), .ZN(n2114) );
  OAI21_X4 U950 ( .B1(n2829), .B2(n3157), .A(n2115), .ZN(n891) );
  AOI222_X2 U951 ( .A1(n3144), .A2(n427), .B1(n333), .B2(n424), .C1(n388), 
        .C2(n421), .ZN(n2115) );
  OAI21_X4 U952 ( .B1(n2830), .B2(n3157), .A(n2116), .ZN(n1734) );
  AOI222_X2 U953 ( .A1(n3145), .A2(n424), .B1(n333), .B2(n421), .C1(n388), 
        .C2(n418), .ZN(n2116) );
  OAI21_X4 U954 ( .B1(n2831), .B2(n3157), .A(n2117), .ZN(n1735) );
  AOI222_X2 U955 ( .A1(n3145), .A2(n421), .B1(n333), .B2(n418), .C1(n388), 
        .C2(n415), .ZN(n2117) );
  OAI21_X4 U956 ( .B1(n2832), .B2(n3157), .A(n2118), .ZN(n1736) );
  AOI222_X2 U957 ( .A1(n3144), .A2(n418), .B1(n333), .B2(n415), .C1(n388), 
        .C2(n412), .ZN(n2118) );
  OAI21_X4 U958 ( .B1(n2833), .B2(n3157), .A(n2119), .ZN(n941) );
  AOI222_X2 U959 ( .A1(n3144), .A2(n415), .B1(n333), .B2(n412), .C1(n388), 
        .C2(n409), .ZN(n2119) );
  OAI21_X4 U960 ( .B1(n2834), .B2(n3156), .A(n2120), .ZN(n1737) );
  AOI222_X2 U961 ( .A1(n3144), .A2(n412), .B1(n333), .B2(n409), .C1(n388), 
        .C2(n406), .ZN(n2120) );
  OAI21_X4 U962 ( .B1(n2835), .B2(n3156), .A(n2121), .ZN(n1738) );
  AOI222_X2 U963 ( .A1(n3145), .A2(n409), .B1(n333), .B2(n406), .C1(n388), 
        .C2(n403), .ZN(n2121) );
  OAI21_X4 U964 ( .B1(n2836), .B2(n3156), .A(n2122), .ZN(n1739) );
  AOI222_X2 U965 ( .A1(n3145), .A2(n406), .B1(n333), .B2(n403), .C1(n388), 
        .C2(n400), .ZN(n2122) );
  OAI21_X4 U966 ( .B1(n2837), .B2(n3156), .A(n2123), .ZN(n1740) );
  AOI222_X2 U967 ( .A1(n3144), .A2(n403), .B1(n333), .B2(n400), .C1(n388), 
        .C2(n397), .ZN(n2123) );
  OAI21_X4 U968 ( .B1(n2838), .B2(n3156), .A(n2124), .ZN(n1741) );
  AOI222_X2 U969 ( .A1(n3145), .A2(n400), .B1(n333), .B2(n397), .C1(n388), 
        .C2(n393), .ZN(n2124) );
  OAI21_X4 U970 ( .B1(n2839), .B2(n3156), .A(n2125), .ZN(n1742) );
  AOI222_X2 U971 ( .A1(n3145), .A2(n397), .B1(n333), .B2(n393), .C1(n388), 
        .C2(n390), .ZN(n2125) );
  OAI21_X4 U972 ( .B1(n2840), .B2(n3156), .A(n2126), .ZN(n1743) );
  OAI21_X4 U974 ( .B1(n2841), .B2(n3156), .A(n2127), .ZN(n1744) );
  AND2_X4 U976 ( .A1(n3144), .A2(n390), .ZN(n1376) );
  XOR2_X2 U978 ( .A(n2128), .B(n289), .Z(n1746) );
  OAI21_X4 U979 ( .B1(n2808), .B2(n3160), .A(n2162), .ZN(n2128) );
  NAND2_X4 U980 ( .A1(n386), .A2(n484), .ZN(n2162) );
  XOR2_X2 U981 ( .A(n2129), .B(n289), .Z(n1747) );
  OAI21_X4 U982 ( .B1(n2809), .B2(n3160), .A(n2163), .ZN(n2129) );
  AOI21_X4 U983 ( .B1(n386), .B2(n481), .A(n1377), .ZN(n2163) );
  AND2_X4 U984 ( .A1(n331), .A2(n484), .ZN(n1377) );
  XOR2_X2 U985 ( .A(n2130), .B(n289), .Z(n1748) );
  OAI21_X4 U986 ( .B1(n2810), .B2(n3160), .A(n2164), .ZN(n2130) );
  AOI222_X2 U987 ( .A1(n3148), .A2(n484), .B1(n331), .B2(n481), .C1(n386), 
        .C2(n478), .ZN(n2164) );
  XOR2_X2 U988 ( .A(n2131), .B(n289), .Z(n1749) );
  OAI21_X4 U989 ( .B1(n2811), .B2(n3160), .A(n2165), .ZN(n2131) );
  AOI222_X2 U990 ( .A1(n3147), .A2(n481), .B1(n331), .B2(n478), .C1(n386), 
        .C2(n475), .ZN(n2165) );
  XOR2_X2 U991 ( .A(n2132), .B(n289), .Z(n1750) );
  OAI21_X4 U992 ( .B1(n2812), .B2(n3160), .A(n2166), .ZN(n2132) );
  AOI222_X2 U993 ( .A1(n3148), .A2(n478), .B1(n331), .B2(n475), .C1(n386), 
        .C2(n472), .ZN(n2166) );
  XOR2_X2 U994 ( .A(n2133), .B(n289), .Z(n1751) );
  OAI21_X4 U995 ( .B1(n2813), .B2(n3160), .A(n2167), .ZN(n2133) );
  AOI222_X2 U996 ( .A1(n3147), .A2(n475), .B1(n331), .B2(n472), .C1(n386), 
        .C2(n469), .ZN(n2167) );
  XOR2_X2 U997 ( .A(n2134), .B(n289), .Z(n1752) );
  OAI21_X4 U998 ( .B1(n2814), .B2(n3160), .A(n2168), .ZN(n2134) );
  AOI222_X2 U999 ( .A1(n3148), .A2(n472), .B1(n331), .B2(n469), .C1(n386), 
        .C2(n466), .ZN(n2168) );
  XOR2_X2 U1000 ( .A(n2135), .B(n289), .Z(n1753) );
  OAI21_X4 U1001 ( .B1(n2815), .B2(n3160), .A(n2169), .ZN(n2135) );
  AOI222_X2 U1002 ( .A1(n3147), .A2(n469), .B1(n331), .B2(n466), .C1(n386), 
        .C2(n463), .ZN(n2169) );
  XOR2_X2 U1003 ( .A(n2136), .B(n289), .Z(n1754) );
  OAI21_X4 U1004 ( .B1(n2816), .B2(n3160), .A(n2170), .ZN(n2136) );
  AOI222_X2 U1005 ( .A1(n3148), .A2(n466), .B1(n331), .B2(n463), .C1(n386), 
        .C2(n460), .ZN(n2170) );
  XOR2_X2 U1006 ( .A(n2137), .B(n289), .Z(n1755) );
  OAI21_X4 U1007 ( .B1(n2817), .B2(n3160), .A(n2171), .ZN(n2137) );
  AOI222_X2 U1008 ( .A1(n3147), .A2(n463), .B1(n331), .B2(n460), .C1(n386), 
        .C2(n457), .ZN(n2171) );
  XOR2_X2 U1009 ( .A(n2138), .B(n289), .Z(n1756) );
  OAI21_X4 U1010 ( .B1(n2818), .B2(n3160), .A(n2172), .ZN(n2138) );
  AOI222_X2 U1011 ( .A1(n3148), .A2(n460), .B1(n331), .B2(n457), .C1(n386), 
        .C2(n454), .ZN(n2172) );
  XOR2_X2 U1012 ( .A(n2139), .B(n289), .Z(n1757) );
  OAI21_X4 U1013 ( .B1(n2819), .B2(n3160), .A(n2173), .ZN(n2139) );
  AOI222_X2 U1014 ( .A1(n3147), .A2(n457), .B1(n331), .B2(n454), .C1(n386), 
        .C2(n451), .ZN(n2173) );
  XOR2_X2 U1015 ( .A(n2140), .B(n289), .Z(n1758) );
  OAI21_X4 U1016 ( .B1(n2820), .B2(n3160), .A(n2174), .ZN(n2140) );
  AOI222_X2 U1017 ( .A1(n3147), .A2(n454), .B1(n331), .B2(n451), .C1(n386), 
        .C2(n448), .ZN(n2174) );
  XOR2_X2 U1018 ( .A(n2141), .B(n289), .Z(n1759) );
  OAI21_X4 U1019 ( .B1(n2821), .B2(n3160), .A(n2175), .ZN(n2141) );
  AOI222_X2 U1020 ( .A1(n3148), .A2(n451), .B1(n331), .B2(n448), .C1(n386), 
        .C2(n445), .ZN(n2175) );
  XOR2_X2 U1021 ( .A(n2142), .B(n289), .Z(n1760) );
  OAI21_X4 U1022 ( .B1(n2822), .B2(n3160), .A(n2176), .ZN(n2142) );
  AOI222_X2 U1023 ( .A1(n3148), .A2(n448), .B1(n331), .B2(n445), .C1(n386), 
        .C2(n442), .ZN(n2176) );
  XOR2_X2 U1024 ( .A(n2143), .B(n289), .Z(n1761) );
  OAI21_X4 U1025 ( .B1(n2823), .B2(n3160), .A(n2177), .ZN(n2143) );
  AOI222_X2 U1026 ( .A1(n3147), .A2(n445), .B1(n331), .B2(n442), .C1(n386), 
        .C2(n439), .ZN(n2177) );
  XOR2_X2 U1027 ( .A(n2144), .B(n289), .Z(n1762) );
  OAI21_X4 U1028 ( .B1(n2824), .B2(n3160), .A(n2178), .ZN(n2144) );
  AOI222_X2 U1029 ( .A1(n3148), .A2(n442), .B1(n331), .B2(n439), .C1(n386), 
        .C2(n436), .ZN(n2178) );
  XOR2_X2 U1030 ( .A(n2145), .B(n289), .Z(n1763) );
  OAI21_X4 U1031 ( .B1(n2825), .B2(n3160), .A(n2179), .ZN(n2145) );
  AOI222_X2 U1032 ( .A1(n3147), .A2(n439), .B1(n331), .B2(n436), .C1(n386), 
        .C2(n433), .ZN(n2179) );
  XOR2_X2 U1033 ( .A(n2146), .B(n289), .Z(n1764) );
  OAI21_X4 U1034 ( .B1(n2826), .B2(n3160), .A(n2180), .ZN(n2146) );
  AOI222_X2 U1035 ( .A1(n3148), .A2(n436), .B1(n331), .B2(n433), .C1(n386), 
        .C2(n430), .ZN(n2180) );
  XOR2_X2 U1036 ( .A(n2147), .B(n289), .Z(n907) );
  OAI21_X4 U1037 ( .B1(n2827), .B2(n3160), .A(n2181), .ZN(n2147) );
  AOI222_X2 U1038 ( .A1(n3147), .A2(n433), .B1(n331), .B2(n430), .C1(n386), 
        .C2(n427), .ZN(n2181) );
  XOR2_X2 U1039 ( .A(n2148), .B(n289), .Z(n1765) );
  OAI21_X4 U1040 ( .B1(n2828), .B2(n3160), .A(n2182), .ZN(n2148) );
  AOI222_X2 U1041 ( .A1(n3148), .A2(n430), .B1(n331), .B2(n427), .C1(n386), 
        .C2(n424), .ZN(n2182) );
  XOR2_X2 U1042 ( .A(n2149), .B(n289), .Z(n1766) );
  OAI21_X4 U1043 ( .B1(n2829), .B2(n3160), .A(n2183), .ZN(n2149) );
  AOI222_X2 U1044 ( .A1(n3147), .A2(n427), .B1(n331), .B2(n424), .C1(n386), 
        .C2(n421), .ZN(n2183) );
  XOR2_X2 U1045 ( .A(n2150), .B(n289), .Z(n1767) );
  OAI21_X4 U1046 ( .B1(n2830), .B2(n3160), .A(n2184), .ZN(n2150) );
  AOI222_X2 U1047 ( .A1(n3148), .A2(n424), .B1(n331), .B2(n421), .C1(n386), 
        .C2(n418), .ZN(n2184) );
  XOR2_X2 U1048 ( .A(n2151), .B(n289), .Z(n1768) );
  OAI21_X4 U1049 ( .B1(n2831), .B2(n3160), .A(n2185), .ZN(n2151) );
  AOI222_X2 U1050 ( .A1(n3147), .A2(n421), .B1(n331), .B2(n418), .C1(n386), 
        .C2(n415), .ZN(n2185) );
  XOR2_X2 U1051 ( .A(n2152), .B(n289), .Z(n1769) );
  OAI21_X4 U1052 ( .B1(n2832), .B2(n3160), .A(n2186), .ZN(n2152) );
  AOI222_X2 U1053 ( .A1(n3148), .A2(n418), .B1(n331), .B2(n415), .C1(n386), 
        .C2(n412), .ZN(n2186) );
  XOR2_X2 U1054 ( .A(n2153), .B(n289), .Z(n1770) );
  OAI21_X4 U1055 ( .B1(n2833), .B2(n3160), .A(n2187), .ZN(n2153) );
  AOI222_X2 U1056 ( .A1(n3147), .A2(n415), .B1(n331), .B2(n412), .C1(n386), 
        .C2(n409), .ZN(n2187) );
  XOR2_X2 U1057 ( .A(n2154), .B(n289), .Z(n1771) );
  OAI21_X4 U1058 ( .B1(n2834), .B2(n3159), .A(n2188), .ZN(n2154) );
  AOI222_X2 U1059 ( .A1(n3148), .A2(n412), .B1(n331), .B2(n409), .C1(n386), 
        .C2(n406), .ZN(n2188) );
  XOR2_X2 U1060 ( .A(n2155), .B(n289), .Z(n1772) );
  OAI21_X4 U1061 ( .B1(n2835), .B2(n3159), .A(n2189), .ZN(n2155) );
  AOI222_X2 U1062 ( .A1(n3147), .A2(n409), .B1(n331), .B2(n406), .C1(n386), 
        .C2(n403), .ZN(n2189) );
  XOR2_X2 U1063 ( .A(n2156), .B(n289), .Z(n1773) );
  OAI21_X4 U1064 ( .B1(n2836), .B2(n3159), .A(n2190), .ZN(n2156) );
  AOI222_X2 U1065 ( .A1(n3148), .A2(n406), .B1(n331), .B2(n403), .C1(n386), 
        .C2(n400), .ZN(n2190) );
  XOR2_X2 U1066 ( .A(n2157), .B(n289), .Z(n1774) );
  OAI21_X4 U1067 ( .B1(n2837), .B2(n3159), .A(n2191), .ZN(n2157) );
  AOI222_X2 U1068 ( .A1(n3147), .A2(n403), .B1(n331), .B2(n400), .C1(n386), 
        .C2(n397), .ZN(n2191) );
  XOR2_X2 U1069 ( .A(n2158), .B(n289), .Z(n1775) );
  OAI21_X4 U1070 ( .B1(n2838), .B2(n3159), .A(n2192), .ZN(n2158) );
  AOI222_X2 U1071 ( .A1(n3148), .A2(n400), .B1(n331), .B2(n397), .C1(n386), 
        .C2(n393), .ZN(n2192) );
  XOR2_X2 U1072 ( .A(n2159), .B(n289), .Z(n1776) );
  OAI21_X4 U1073 ( .B1(n2839), .B2(n3159), .A(n2193), .ZN(n2159) );
  AOI222_X2 U1074 ( .A1(n3147), .A2(n397), .B1(n331), .B2(n393), .C1(n386), 
        .C2(n390), .ZN(n2193) );
  XOR2_X2 U1075 ( .A(n2160), .B(n289), .Z(n1777) );
  OAI21_X4 U1076 ( .B1(n2840), .B2(n3159), .A(n2194), .ZN(n2160) );
  XOR2_X2 U1078 ( .A(n2161), .B(n289), .Z(n1778) );
  OAI21_X4 U1079 ( .B1(n2841), .B2(n3159), .A(n2195), .ZN(n2161) );
  AND2_X4 U1081 ( .A1(n3147), .A2(n390), .ZN(n1379) );
  XOR2_X2 U1083 ( .A(n2196), .B(n286), .Z(n1780) );
  OAI21_X4 U1084 ( .B1(n2808), .B2(n3161), .A(n2230), .ZN(n2196) );
  NAND2_X4 U1085 ( .A1(n384), .A2(n484), .ZN(n2230) );
  XOR2_X2 U1086 ( .A(n2197), .B(n286), .Z(n1781) );
  OAI21_X4 U1087 ( .B1(n2809), .B2(n3161), .A(n2231), .ZN(n2197) );
  AOI21_X4 U1088 ( .B1(n384), .B2(n481), .A(n1380), .ZN(n2231) );
  AND2_X4 U1089 ( .A1(n329), .A2(n484), .ZN(n1380) );
  XOR2_X2 U1090 ( .A(n2198), .B(n286), .Z(n1782) );
  OAI21_X4 U1091 ( .B1(n2810), .B2(n360), .A(n2232), .ZN(n2198) );
  AOI222_X2 U1092 ( .A1(n3151), .A2(n484), .B1(n329), .B2(n481), .C1(n384), 
        .C2(n478), .ZN(n2232) );
  XOR2_X2 U1093 ( .A(n2199), .B(n286), .Z(n1783) );
  OAI21_X4 U1094 ( .B1(n2811), .B2(n360), .A(n2233), .ZN(n2199) );
  AOI222_X2 U1095 ( .A1(n3150), .A2(n481), .B1(n329), .B2(n478), .C1(n384), 
        .C2(n475), .ZN(n2233) );
  XOR2_X2 U1096 ( .A(n2200), .B(n286), .Z(n1784) );
  OAI21_X4 U1097 ( .B1(n2812), .B2(n360), .A(n2234), .ZN(n2200) );
  AOI222_X2 U1098 ( .A1(n3151), .A2(n478), .B1(n329), .B2(n475), .C1(n384), 
        .C2(n472), .ZN(n2234) );
  XOR2_X2 U1099 ( .A(n2201), .B(n286), .Z(n1785) );
  OAI21_X4 U1100 ( .B1(n2813), .B2(n360), .A(n2235), .ZN(n2201) );
  AOI222_X2 U1101 ( .A1(n3150), .A2(n475), .B1(n329), .B2(n472), .C1(n384), 
        .C2(n469), .ZN(n2235) );
  XOR2_X2 U1102 ( .A(n2202), .B(n286), .Z(n1786) );
  OAI21_X4 U1103 ( .B1(n2814), .B2(n360), .A(n2236), .ZN(n2202) );
  AOI222_X2 U1104 ( .A1(n3151), .A2(n472), .B1(n329), .B2(n469), .C1(n384), 
        .C2(n466), .ZN(n2236) );
  XOR2_X2 U1105 ( .A(n2203), .B(n286), .Z(n1787) );
  OAI21_X4 U1106 ( .B1(n2815), .B2(n360), .A(n2237), .ZN(n2203) );
  AOI222_X2 U1107 ( .A1(n3150), .A2(n469), .B1(n329), .B2(n466), .C1(n384), 
        .C2(n463), .ZN(n2237) );
  XOR2_X2 U1108 ( .A(n2204), .B(n286), .Z(n1788) );
  OAI21_X4 U1109 ( .B1(n2816), .B2(n360), .A(n2238), .ZN(n2204) );
  AOI222_X2 U1110 ( .A1(n3151), .A2(n466), .B1(n329), .B2(n463), .C1(n384), 
        .C2(n460), .ZN(n2238) );
  XOR2_X2 U1111 ( .A(n2205), .B(n286), .Z(n1789) );
  OAI21_X4 U1112 ( .B1(n2817), .B2(n360), .A(n2239), .ZN(n2205) );
  AOI222_X2 U1113 ( .A1(n3150), .A2(n463), .B1(n329), .B2(n460), .C1(n384), 
        .C2(n457), .ZN(n2239) );
  XOR2_X2 U1114 ( .A(n2206), .B(n286), .Z(n1790) );
  OAI21_X4 U1115 ( .B1(n2818), .B2(n360), .A(n2240), .ZN(n2206) );
  AOI222_X2 U1116 ( .A1(n3151), .A2(n460), .B1(n329), .B2(n457), .C1(n384), 
        .C2(n454), .ZN(n2240) );
  XOR2_X2 U1117 ( .A(n2207), .B(n286), .Z(n1791) );
  OAI21_X4 U1118 ( .B1(n2819), .B2(n360), .A(n2241), .ZN(n2207) );
  AOI222_X2 U1119 ( .A1(n3150), .A2(n457), .B1(n329), .B2(n454), .C1(n384), 
        .C2(n451), .ZN(n2241) );
  XOR2_X2 U1120 ( .A(n2208), .B(n286), .Z(n1792) );
  OAI21_X4 U1121 ( .B1(n2820), .B2(n360), .A(n2242), .ZN(n2208) );
  AOI222_X2 U1122 ( .A1(n3151), .A2(n454), .B1(n329), .B2(n451), .C1(n384), 
        .C2(n448), .ZN(n2242) );
  XOR2_X2 U1123 ( .A(n2209), .B(n286), .Z(n1793) );
  OAI21_X4 U1124 ( .B1(n2821), .B2(n360), .A(n2243), .ZN(n2209) );
  AOI222_X2 U1125 ( .A1(n3150), .A2(n451), .B1(n329), .B2(n448), .C1(n384), 
        .C2(n445), .ZN(n2243) );
  XOR2_X2 U1126 ( .A(n2210), .B(n286), .Z(n1794) );
  OAI21_X4 U1127 ( .B1(n2822), .B2(n360), .A(n2244), .ZN(n2210) );
  AOI222_X2 U1128 ( .A1(n3151), .A2(n448), .B1(n329), .B2(n445), .C1(n384), 
        .C2(n442), .ZN(n2244) );
  XOR2_X2 U1129 ( .A(n2211), .B(n286), .Z(n1795) );
  OAI21_X4 U1130 ( .B1(n2823), .B2(n360), .A(n2245), .ZN(n2211) );
  AOI222_X2 U1131 ( .A1(n3150), .A2(n445), .B1(n329), .B2(n442), .C1(n384), 
        .C2(n439), .ZN(n2245) );
  XOR2_X2 U1132 ( .A(n2212), .B(n286), .Z(n1796) );
  OAI21_X4 U1133 ( .B1(n2824), .B2(n360), .A(n2246), .ZN(n2212) );
  AOI222_X2 U1134 ( .A1(n3151), .A2(n442), .B1(n329), .B2(n439), .C1(n384), 
        .C2(n436), .ZN(n2246) );
  XOR2_X2 U1135 ( .A(n2213), .B(n286), .Z(n1797) );
  OAI21_X4 U1136 ( .B1(n2825), .B2(n360), .A(n2247), .ZN(n2213) );
  AOI222_X2 U1137 ( .A1(n3150), .A2(n439), .B1(n329), .B2(n436), .C1(n384), 
        .C2(n433), .ZN(n2247) );
  XOR2_X2 U1138 ( .A(n2214), .B(n286), .Z(n1798) );
  OAI21_X4 U1139 ( .B1(n2826), .B2(n360), .A(n2248), .ZN(n2214) );
  AOI222_X2 U1140 ( .A1(n3151), .A2(n436), .B1(n329), .B2(n433), .C1(n384), 
        .C2(n430), .ZN(n2248) );
  XOR2_X2 U1141 ( .A(n2215), .B(n286), .Z(n1799) );
  OAI21_X4 U1142 ( .B1(n2827), .B2(n360), .A(n2249), .ZN(n2215) );
  AOI222_X2 U1143 ( .A1(n3150), .A2(n433), .B1(n329), .B2(n430), .C1(n384), 
        .C2(n427), .ZN(n2249) );
  XOR2_X2 U1144 ( .A(n2216), .B(n286), .Z(n1800) );
  OAI21_X4 U1145 ( .B1(n2828), .B2(n360), .A(n2250), .ZN(n2216) );
  AOI222_X2 U1146 ( .A1(n3151), .A2(n430), .B1(n329), .B2(n427), .C1(n384), 
        .C2(n424), .ZN(n2250) );
  XOR2_X2 U1147 ( .A(n2217), .B(n286), .Z(n1801) );
  OAI21_X4 U1148 ( .B1(n2829), .B2(n360), .A(n2251), .ZN(n2217) );
  AOI222_X2 U1149 ( .A1(n3150), .A2(n427), .B1(n329), .B2(n424), .C1(n384), 
        .C2(n421), .ZN(n2251) );
  XOR2_X2 U1150 ( .A(n2218), .B(n286), .Z(n1802) );
  OAI21_X4 U1151 ( .B1(n2830), .B2(n360), .A(n2252), .ZN(n2218) );
  AOI222_X2 U1152 ( .A1(n3151), .A2(n424), .B1(n329), .B2(n421), .C1(n384), 
        .C2(n418), .ZN(n2252) );
  XOR2_X2 U1153 ( .A(n2219), .B(n286), .Z(n1803) );
  OAI21_X4 U1154 ( .B1(n2831), .B2(n360), .A(n2253), .ZN(n2219) );
  AOI222_X2 U1155 ( .A1(n3150), .A2(n421), .B1(n329), .B2(n418), .C1(n384), 
        .C2(n415), .ZN(n2253) );
  XOR2_X2 U1156 ( .A(n2220), .B(n286), .Z(n1804) );
  OAI21_X4 U1157 ( .B1(n2832), .B2(n360), .A(n2254), .ZN(n2220) );
  AOI222_X2 U1158 ( .A1(n3151), .A2(n418), .B1(n329), .B2(n415), .C1(n384), 
        .C2(n412), .ZN(n2254) );
  XOR2_X2 U1159 ( .A(n2221), .B(n286), .Z(n1805) );
  OAI21_X4 U1160 ( .B1(n2833), .B2(n360), .A(n2255), .ZN(n2221) );
  AOI222_X2 U1161 ( .A1(n3150), .A2(n415), .B1(n329), .B2(n412), .C1(n384), 
        .C2(n409), .ZN(n2255) );
  XOR2_X2 U1162 ( .A(n2222), .B(n286), .Z(n1806) );
  OAI21_X4 U1163 ( .B1(n2834), .B2(n360), .A(n2256), .ZN(n2222) );
  AOI222_X2 U1164 ( .A1(n3151), .A2(n412), .B1(n329), .B2(n409), .C1(n384), 
        .C2(n406), .ZN(n2256) );
  XOR2_X2 U1165 ( .A(n2223), .B(n286), .Z(n1807) );
  OAI21_X4 U1166 ( .B1(n2835), .B2(n360), .A(n2257), .ZN(n2223) );
  AOI222_X2 U1167 ( .A1(n3151), .A2(n409), .B1(n329), .B2(n406), .C1(n384), 
        .C2(n403), .ZN(n2257) );
  XOR2_X2 U1168 ( .A(n2224), .B(n286), .Z(n1808) );
  OAI21_X4 U1169 ( .B1(n2836), .B2(n360), .A(n2258), .ZN(n2224) );
  AOI222_X2 U1170 ( .A1(n3150), .A2(n406), .B1(n329), .B2(n403), .C1(n384), 
        .C2(n400), .ZN(n2258) );
  XOR2_X2 U1171 ( .A(n2225), .B(n286), .Z(n1809) );
  OAI21_X4 U1172 ( .B1(n2837), .B2(n360), .A(n2259), .ZN(n2225) );
  AOI222_X2 U1173 ( .A1(n3150), .A2(n403), .B1(n329), .B2(n400), .C1(n384), 
        .C2(n397), .ZN(n2259) );
  XOR2_X2 U1174 ( .A(n2226), .B(n286), .Z(n1810) );
  OAI21_X4 U1175 ( .B1(n2838), .B2(n360), .A(n2260), .ZN(n2226) );
  AOI222_X2 U1176 ( .A1(n3151), .A2(n400), .B1(n329), .B2(n397), .C1(n384), 
        .C2(n393), .ZN(n2260) );
  XOR2_X2 U1177 ( .A(n2227), .B(n286), .Z(n1811) );
  OAI21_X4 U1178 ( .B1(n2839), .B2(n360), .A(n2261), .ZN(n2227) );
  AOI222_X2 U1179 ( .A1(n3150), .A2(n397), .B1(n329), .B2(n393), .C1(n384), 
        .C2(n390), .ZN(n2261) );
  XOR2_X2 U1180 ( .A(n2228), .B(n286), .Z(n1812) );
  OAI21_X4 U1181 ( .B1(n2840), .B2(n360), .A(n2262), .ZN(n2228) );
  XOR2_X2 U1183 ( .A(n2229), .B(n286), .Z(n1813) );
  OAI21_X4 U1184 ( .B1(n2841), .B2(n360), .A(n2263), .ZN(n2229) );
  AND2_X4 U1186 ( .A1(n3150), .A2(n390), .ZN(n1382) );
  XOR2_X2 U1188 ( .A(n2264), .B(n283), .Z(n1815) );
  OAI21_X4 U1189 ( .B1(n2808), .B2(n3162), .A(n2298), .ZN(n2264) );
  NAND2_X4 U1190 ( .A1(n382), .A2(n484), .ZN(n2298) );
  XOR2_X2 U1191 ( .A(n2265), .B(n283), .Z(n1816) );
  OAI21_X4 U1192 ( .B1(n2809), .B2(n3162), .A(n2299), .ZN(n2265) );
  AOI21_X4 U1193 ( .B1(n382), .B2(n481), .A(n1383), .ZN(n2299) );
  AND2_X4 U1194 ( .A1(n327), .A2(n484), .ZN(n1383) );
  XOR2_X2 U1195 ( .A(n2266), .B(n283), .Z(n1817) );
  OAI21_X4 U1196 ( .B1(n2810), .B2(n357), .A(n2300), .ZN(n2266) );
  AOI222_X2 U1197 ( .A1(n3136), .A2(n484), .B1(n327), .B2(n481), .C1(n382), 
        .C2(n478), .ZN(n2300) );
  XOR2_X2 U1198 ( .A(n2267), .B(n283), .Z(n1818) );
  OAI21_X4 U1199 ( .B1(n2811), .B2(n357), .A(n2301), .ZN(n2267) );
  AOI222_X2 U1200 ( .A1(n3135), .A2(n481), .B1(n327), .B2(n478), .C1(n382), 
        .C2(n475), .ZN(n2301) );
  XOR2_X2 U1201 ( .A(n2268), .B(n283), .Z(n1819) );
  OAI21_X4 U1202 ( .B1(n2812), .B2(n357), .A(n2302), .ZN(n2268) );
  AOI222_X2 U1203 ( .A1(n3136), .A2(n478), .B1(n327), .B2(n475), .C1(n382), 
        .C2(n472), .ZN(n2302) );
  XOR2_X2 U1204 ( .A(n2269), .B(n283), .Z(n1820) );
  OAI21_X4 U1205 ( .B1(n2813), .B2(n357), .A(n2303), .ZN(n2269) );
  AOI222_X2 U1206 ( .A1(n3135), .A2(n475), .B1(n327), .B2(n472), .C1(n382), 
        .C2(n469), .ZN(n2303) );
  XOR2_X2 U1207 ( .A(n2270), .B(n283), .Z(n1821) );
  OAI21_X4 U1208 ( .B1(n2814), .B2(n357), .A(n2304), .ZN(n2270) );
  AOI222_X2 U1209 ( .A1(n3136), .A2(n472), .B1(n327), .B2(n469), .C1(n382), 
        .C2(n466), .ZN(n2304) );
  XOR2_X2 U1210 ( .A(n2271), .B(n283), .Z(n1822) );
  OAI21_X4 U1211 ( .B1(n2815), .B2(n357), .A(n2305), .ZN(n2271) );
  AOI222_X2 U1212 ( .A1(n3135), .A2(n469), .B1(n327), .B2(n466), .C1(n382), 
        .C2(n463), .ZN(n2305) );
  XOR2_X2 U1213 ( .A(n2272), .B(n283), .Z(n1823) );
  OAI21_X4 U1214 ( .B1(n2816), .B2(n357), .A(n2306), .ZN(n2272) );
  AOI222_X2 U1215 ( .A1(n3136), .A2(n466), .B1(n327), .B2(n463), .C1(n382), 
        .C2(n460), .ZN(n2306) );
  XOR2_X2 U1216 ( .A(n2273), .B(n283), .Z(n1824) );
  OAI21_X4 U1217 ( .B1(n2817), .B2(n357), .A(n2307), .ZN(n2273) );
  AOI222_X2 U1218 ( .A1(n3135), .A2(n463), .B1(n327), .B2(n460), .C1(n382), 
        .C2(n457), .ZN(n2307) );
  XOR2_X2 U1219 ( .A(n2274), .B(n283), .Z(n1825) );
  OAI21_X4 U1220 ( .B1(n2818), .B2(n357), .A(n2308), .ZN(n2274) );
  AOI222_X2 U1221 ( .A1(n3136), .A2(n460), .B1(n327), .B2(n457), .C1(n382), 
        .C2(n454), .ZN(n2308) );
  XOR2_X2 U1222 ( .A(n2275), .B(n283), .Z(n1826) );
  OAI21_X4 U1223 ( .B1(n2819), .B2(n357), .A(n2309), .ZN(n2275) );
  AOI222_X2 U1224 ( .A1(n3135), .A2(n457), .B1(n327), .B2(n454), .C1(n382), 
        .C2(n451), .ZN(n2309) );
  XOR2_X2 U1225 ( .A(n2276), .B(n283), .Z(n1827) );
  OAI21_X4 U1226 ( .B1(n2820), .B2(n357), .A(n2310), .ZN(n2276) );
  AOI222_X2 U1227 ( .A1(n3136), .A2(n454), .B1(n327), .B2(n451), .C1(n382), 
        .C2(n448), .ZN(n2310) );
  XOR2_X2 U1228 ( .A(n2277), .B(n283), .Z(n1828) );
  OAI21_X4 U1229 ( .B1(n2821), .B2(n357), .A(n2311), .ZN(n2277) );
  AOI222_X2 U1230 ( .A1(n3135), .A2(n451), .B1(n327), .B2(n448), .C1(n382), 
        .C2(n445), .ZN(n2311) );
  XOR2_X2 U1231 ( .A(n2278), .B(n283), .Z(n1829) );
  OAI21_X4 U1232 ( .B1(n2822), .B2(n357), .A(n2312), .ZN(n2278) );
  AOI222_X2 U1233 ( .A1(n3136), .A2(n448), .B1(n327), .B2(n445), .C1(n382), 
        .C2(n442), .ZN(n2312) );
  XOR2_X2 U1234 ( .A(n2279), .B(n283), .Z(n1830) );
  OAI21_X4 U1235 ( .B1(n2823), .B2(n357), .A(n2313), .ZN(n2279) );
  AOI222_X2 U1236 ( .A1(n3135), .A2(n445), .B1(n327), .B2(n442), .C1(n382), 
        .C2(n439), .ZN(n2313) );
  XOR2_X2 U1237 ( .A(n2280), .B(n283), .Z(n1831) );
  OAI21_X4 U1238 ( .B1(n2824), .B2(n357), .A(n2314), .ZN(n2280) );
  AOI222_X2 U1239 ( .A1(n3136), .A2(n442), .B1(n327), .B2(n439), .C1(n382), 
        .C2(n436), .ZN(n2314) );
  XOR2_X2 U1240 ( .A(n2281), .B(n283), .Z(n1832) );
  OAI21_X4 U1241 ( .B1(n2825), .B2(n357), .A(n2315), .ZN(n2281) );
  AOI222_X2 U1242 ( .A1(n3135), .A2(n439), .B1(n327), .B2(n436), .C1(n382), 
        .C2(n433), .ZN(n2315) );
  XOR2_X2 U1243 ( .A(n2282), .B(n283), .Z(n1833) );
  OAI21_X4 U1244 ( .B1(n2826), .B2(n357), .A(n2316), .ZN(n2282) );
  AOI222_X2 U1245 ( .A1(n3136), .A2(n436), .B1(n327), .B2(n433), .C1(n382), 
        .C2(n430), .ZN(n2316) );
  XOR2_X2 U1246 ( .A(n2283), .B(n283), .Z(n1834) );
  OAI21_X4 U1247 ( .B1(n2827), .B2(n357), .A(n2317), .ZN(n2283) );
  AOI222_X2 U1248 ( .A1(n3135), .A2(n433), .B1(n327), .B2(n430), .C1(n382), 
        .C2(n427), .ZN(n2317) );
  XOR2_X2 U1249 ( .A(n2284), .B(n283), .Z(n1835) );
  OAI21_X4 U1250 ( .B1(n2828), .B2(n357), .A(n2318), .ZN(n2284) );
  AOI222_X2 U1251 ( .A1(n3136), .A2(n430), .B1(n327), .B2(n427), .C1(n382), 
        .C2(n424), .ZN(n2318) );
  XOR2_X2 U1252 ( .A(n2285), .B(n283), .Z(n1836) );
  OAI21_X4 U1253 ( .B1(n2829), .B2(n357), .A(n2319), .ZN(n2285) );
  AOI222_X2 U1254 ( .A1(n3136), .A2(n427), .B1(n327), .B2(n424), .C1(n382), 
        .C2(n421), .ZN(n2319) );
  XOR2_X2 U1255 ( .A(n2286), .B(n283), .Z(n1837) );
  OAI21_X4 U1256 ( .B1(n2830), .B2(n357), .A(n2320), .ZN(n2286) );
  AOI222_X2 U1257 ( .A1(n3135), .A2(n424), .B1(n327), .B2(n421), .C1(n382), 
        .C2(n418), .ZN(n2320) );
  XOR2_X2 U1258 ( .A(n2287), .B(n283), .Z(n1838) );
  OAI21_X4 U1259 ( .B1(n2831), .B2(n357), .A(n2321), .ZN(n2287) );
  AOI222_X2 U1260 ( .A1(n3135), .A2(n421), .B1(n327), .B2(n418), .C1(n382), 
        .C2(n415), .ZN(n2321) );
  XOR2_X2 U1261 ( .A(n2288), .B(n283), .Z(n1839) );
  OAI21_X4 U1262 ( .B1(n2832), .B2(n357), .A(n2322), .ZN(n2288) );
  AOI222_X2 U1263 ( .A1(n3135), .A2(n418), .B1(n327), .B2(n415), .C1(n382), 
        .C2(n412), .ZN(n2322) );
  XOR2_X2 U1264 ( .A(n2289), .B(n283), .Z(n1840) );
  OAI21_X4 U1265 ( .B1(n2833), .B2(n357), .A(n2323), .ZN(n2289) );
  AOI222_X2 U1266 ( .A1(n3136), .A2(n415), .B1(n327), .B2(n412), .C1(n382), 
        .C2(n409), .ZN(n2323) );
  XOR2_X2 U1267 ( .A(n2290), .B(n283), .Z(n1841) );
  OAI21_X4 U1268 ( .B1(n2834), .B2(n357), .A(n2324), .ZN(n2290) );
  AOI222_X2 U1269 ( .A1(n3136), .A2(n412), .B1(n327), .B2(n409), .C1(n382), 
        .C2(n406), .ZN(n2324) );
  XOR2_X2 U1270 ( .A(n2291), .B(n283), .Z(n1842) );
  OAI21_X4 U1271 ( .B1(n2835), .B2(n357), .A(n2325), .ZN(n2291) );
  AOI222_X2 U1272 ( .A1(n3136), .A2(n409), .B1(n327), .B2(n406), .C1(n382), 
        .C2(n403), .ZN(n2325) );
  XOR2_X2 U1273 ( .A(n2292), .B(n283), .Z(n1843) );
  OAI21_X4 U1274 ( .B1(n2836), .B2(n357), .A(n2326), .ZN(n2292) );
  AOI222_X2 U1275 ( .A1(n3135), .A2(n406), .B1(n327), .B2(n403), .C1(n382), 
        .C2(n400), .ZN(n2326) );
  XOR2_X2 U1276 ( .A(n2293), .B(n283), .Z(n1844) );
  OAI21_X4 U1277 ( .B1(n2837), .B2(n357), .A(n2327), .ZN(n2293) );
  AOI222_X2 U1278 ( .A1(n3135), .A2(n403), .B1(n327), .B2(n400), .C1(n382), 
        .C2(n397), .ZN(n2327) );
  XOR2_X2 U1279 ( .A(n2294), .B(n283), .Z(n1845) );
  OAI21_X4 U1280 ( .B1(n2838), .B2(n357), .A(n2328), .ZN(n2294) );
  AOI222_X2 U1281 ( .A1(n3136), .A2(n400), .B1(n327), .B2(n397), .C1(n382), 
        .C2(n393), .ZN(n2328) );
  XOR2_X2 U1282 ( .A(n2295), .B(n283), .Z(n1846) );
  OAI21_X4 U1283 ( .B1(n2839), .B2(n357), .A(n2329), .ZN(n2295) );
  AOI222_X2 U1284 ( .A1(n3135), .A2(n397), .B1(n327), .B2(n393), .C1(n382), 
        .C2(n390), .ZN(n2329) );
  XOR2_X2 U1285 ( .A(n2296), .B(n283), .Z(n1847) );
  OAI21_X4 U1286 ( .B1(n2840), .B2(n357), .A(n2330), .ZN(n2296) );
  XOR2_X2 U1288 ( .A(n2297), .B(n283), .Z(n1848) );
  OAI21_X4 U1289 ( .B1(n2841), .B2(n357), .A(n2331), .ZN(n2297) );
  AND2_X4 U1291 ( .A1(n3135), .A2(n390), .ZN(n1385) );
  XOR2_X2 U1293 ( .A(n2332), .B(n280), .Z(n1850) );
  OAI21_X4 U1294 ( .B1(n2808), .B2(n3129), .A(n2366), .ZN(n2332) );
  NAND2_X4 U1295 ( .A1(n380), .A2(n484), .ZN(n2366) );
  XOR2_X2 U1296 ( .A(n2333), .B(n280), .Z(n1851) );
  OAI21_X4 U1297 ( .B1(n2809), .B2(n3129), .A(n2367), .ZN(n2333) );
  AOI21_X4 U1298 ( .B1(n380), .B2(n481), .A(n1386), .ZN(n2367) );
  AND2_X4 U1299 ( .A1(n325), .A2(n484), .ZN(n1386) );
  XOR2_X2 U1300 ( .A(n2334), .B(n280), .Z(n1852) );
  OAI21_X4 U1301 ( .B1(n2810), .B2(n354), .A(n2368), .ZN(n2334) );
  AOI222_X2 U1302 ( .A1(n3139), .A2(n484), .B1(n325), .B2(n481), .C1(n380), 
        .C2(n478), .ZN(n2368) );
  XOR2_X2 U1303 ( .A(n2335), .B(n280), .Z(n1853) );
  OAI21_X4 U1304 ( .B1(n2811), .B2(n354), .A(n2369), .ZN(n2335) );
  AOI222_X2 U1305 ( .A1(n3138), .A2(n481), .B1(n325), .B2(n478), .C1(n380), 
        .C2(n475), .ZN(n2369) );
  XOR2_X2 U1306 ( .A(n2336), .B(n280), .Z(n1854) );
  OAI21_X4 U1307 ( .B1(n2812), .B2(n354), .A(n2370), .ZN(n2336) );
  AOI222_X2 U1308 ( .A1(n3139), .A2(n478), .B1(n325), .B2(n475), .C1(n380), 
        .C2(n472), .ZN(n2370) );
  XOR2_X2 U1309 ( .A(n2337), .B(n280), .Z(n1855) );
  OAI21_X4 U1310 ( .B1(n2813), .B2(n354), .A(n2371), .ZN(n2337) );
  AOI222_X2 U1311 ( .A1(n3138), .A2(n475), .B1(n325), .B2(n472), .C1(n380), 
        .C2(n469), .ZN(n2371) );
  XOR2_X2 U1312 ( .A(n2338), .B(n280), .Z(n1856) );
  OAI21_X4 U1313 ( .B1(n2814), .B2(n354), .A(n2372), .ZN(n2338) );
  AOI222_X2 U1314 ( .A1(n3139), .A2(n472), .B1(n325), .B2(n469), .C1(n380), 
        .C2(n466), .ZN(n2372) );
  XOR2_X2 U1315 ( .A(n2339), .B(n280), .Z(n1857) );
  OAI21_X4 U1316 ( .B1(n2815), .B2(n354), .A(n2373), .ZN(n2339) );
  AOI222_X2 U1317 ( .A1(n3138), .A2(n469), .B1(n325), .B2(n466), .C1(n380), 
        .C2(n463), .ZN(n2373) );
  XOR2_X2 U1318 ( .A(n2340), .B(n280), .Z(n1858) );
  OAI21_X4 U1319 ( .B1(n2816), .B2(n354), .A(n2374), .ZN(n2340) );
  AOI222_X2 U1320 ( .A1(n3139), .A2(n466), .B1(n325), .B2(n463), .C1(n380), 
        .C2(n460), .ZN(n2374) );
  XOR2_X2 U1321 ( .A(n2341), .B(n280), .Z(n1859) );
  OAI21_X4 U1322 ( .B1(n2817), .B2(n354), .A(n2375), .ZN(n2341) );
  AOI222_X2 U1323 ( .A1(n3138), .A2(n463), .B1(n325), .B2(n460), .C1(n380), 
        .C2(n457), .ZN(n2375) );
  XOR2_X2 U1324 ( .A(n2342), .B(n280), .Z(n1860) );
  OAI21_X4 U1325 ( .B1(n2818), .B2(n354), .A(n2376), .ZN(n2342) );
  AOI222_X2 U1326 ( .A1(n3139), .A2(n460), .B1(n325), .B2(n457), .C1(n380), 
        .C2(n454), .ZN(n2376) );
  XOR2_X2 U1327 ( .A(n2343), .B(n280), .Z(n1861) );
  OAI21_X4 U1328 ( .B1(n2819), .B2(n354), .A(n2377), .ZN(n2343) );
  AOI222_X2 U1329 ( .A1(n3138), .A2(n457), .B1(n325), .B2(n454), .C1(n380), 
        .C2(n451), .ZN(n2377) );
  XOR2_X2 U1330 ( .A(n2344), .B(n280), .Z(n1862) );
  OAI21_X4 U1331 ( .B1(n2820), .B2(n354), .A(n2378), .ZN(n2344) );
  AOI222_X2 U1332 ( .A1(n3139), .A2(n454), .B1(n325), .B2(n451), .C1(n380), 
        .C2(n448), .ZN(n2378) );
  XOR2_X2 U1333 ( .A(n2345), .B(n280), .Z(n1863) );
  OAI21_X4 U1334 ( .B1(n2821), .B2(n354), .A(n2379), .ZN(n2345) );
  AOI222_X2 U1335 ( .A1(n3138), .A2(n451), .B1(n325), .B2(n448), .C1(n380), 
        .C2(n445), .ZN(n2379) );
  XOR2_X2 U1336 ( .A(n2346), .B(n280), .Z(n1864) );
  OAI21_X4 U1337 ( .B1(n2822), .B2(n354), .A(n2380), .ZN(n2346) );
  AOI222_X2 U1338 ( .A1(n3138), .A2(n448), .B1(n325), .B2(n445), .C1(n380), 
        .C2(n442), .ZN(n2380) );
  XOR2_X2 U1339 ( .A(n2347), .B(n280), .Z(n1865) );
  OAI21_X4 U1340 ( .B1(n2823), .B2(n354), .A(n2381), .ZN(n2347) );
  AOI222_X2 U1341 ( .A1(n3139), .A2(n445), .B1(n325), .B2(n442), .C1(n380), 
        .C2(n439), .ZN(n2381) );
  XOR2_X2 U1342 ( .A(n2348), .B(n280), .Z(n1866) );
  OAI21_X4 U1343 ( .B1(n2824), .B2(n354), .A(n2382), .ZN(n2348) );
  AOI222_X2 U1344 ( .A1(n3139), .A2(n442), .B1(n325), .B2(n439), .C1(n380), 
        .C2(n436), .ZN(n2382) );
  XOR2_X2 U1345 ( .A(n2349), .B(n280), .Z(n1867) );
  OAI21_X4 U1346 ( .B1(n2825), .B2(n354), .A(n2383), .ZN(n2349) );
  AOI222_X2 U1347 ( .A1(n3138), .A2(n439), .B1(n325), .B2(n436), .C1(n380), 
        .C2(n433), .ZN(n2383) );
  XOR2_X2 U1348 ( .A(n2350), .B(n280), .Z(n1868) );
  OAI21_X4 U1349 ( .B1(n2826), .B2(n354), .A(n2384), .ZN(n2350) );
  AOI222_X2 U1350 ( .A1(n3139), .A2(n436), .B1(n325), .B2(n433), .C1(n380), 
        .C2(n430), .ZN(n2384) );
  XOR2_X2 U1351 ( .A(n2351), .B(n280), .Z(n1869) );
  OAI21_X4 U1352 ( .B1(n2827), .B2(n354), .A(n2385), .ZN(n2351) );
  AOI222_X2 U1353 ( .A1(n3138), .A2(n433), .B1(n325), .B2(n430), .C1(n380), 
        .C2(n427), .ZN(n2385) );
  XOR2_X2 U1354 ( .A(n2352), .B(n280), .Z(n1870) );
  OAI21_X4 U1355 ( .B1(n2828), .B2(n354), .A(n2386), .ZN(n2352) );
  AOI222_X2 U1356 ( .A1(n3138), .A2(n430), .B1(n325), .B2(n427), .C1(n380), 
        .C2(n424), .ZN(n2386) );
  XOR2_X2 U1357 ( .A(n2353), .B(n280), .Z(n1871) );
  OAI21_X4 U1358 ( .B1(n2829), .B2(n354), .A(n2387), .ZN(n2353) );
  AOI222_X2 U1359 ( .A1(n3139), .A2(n427), .B1(n325), .B2(n424), .C1(n380), 
        .C2(n421), .ZN(n2387) );
  XOR2_X2 U1360 ( .A(n2354), .B(n280), .Z(n1872) );
  OAI21_X4 U1361 ( .B1(n2830), .B2(n354), .A(n2388), .ZN(n2354) );
  AOI222_X2 U1362 ( .A1(n3139), .A2(n424), .B1(n325), .B2(n421), .C1(n380), 
        .C2(n418), .ZN(n2388) );
  XOR2_X2 U1363 ( .A(n2355), .B(n280), .Z(n1873) );
  OAI21_X4 U1364 ( .B1(n2831), .B2(n354), .A(n2389), .ZN(n2355) );
  AOI222_X2 U1365 ( .A1(n3138), .A2(n421), .B1(n325), .B2(n418), .C1(n380), 
        .C2(n415), .ZN(n2389) );
  XOR2_X2 U1366 ( .A(n2356), .B(n280), .Z(n1874) );
  OAI21_X4 U1367 ( .B1(n2832), .B2(n354), .A(n2390), .ZN(n2356) );
  AOI222_X2 U1368 ( .A1(n3138), .A2(n418), .B1(n325), .B2(n415), .C1(n380), 
        .C2(n412), .ZN(n2390) );
  XOR2_X2 U1369 ( .A(n2357), .B(n280), .Z(n1875) );
  OAI21_X4 U1370 ( .B1(n2833), .B2(n354), .A(n2391), .ZN(n2357) );
  AOI222_X2 U1371 ( .A1(n3139), .A2(n415), .B1(n325), .B2(n412), .C1(n380), 
        .C2(n409), .ZN(n2391) );
  XOR2_X2 U1372 ( .A(n2358), .B(n280), .Z(n1876) );
  OAI21_X4 U1373 ( .B1(n2834), .B2(n354), .A(n2392), .ZN(n2358) );
  AOI222_X2 U1374 ( .A1(n3139), .A2(n412), .B1(n325), .B2(n409), .C1(n380), 
        .C2(n406), .ZN(n2392) );
  XOR2_X2 U1375 ( .A(n2359), .B(n280), .Z(n1877) );
  OAI21_X4 U1376 ( .B1(n2835), .B2(n354), .A(n2393), .ZN(n2359) );
  AOI222_X2 U1377 ( .A1(n3139), .A2(n409), .B1(n325), .B2(n406), .C1(n380), 
        .C2(n403), .ZN(n2393) );
  XOR2_X2 U1378 ( .A(n2360), .B(n280), .Z(n1878) );
  OAI21_X4 U1379 ( .B1(n2836), .B2(n354), .A(n2394), .ZN(n2360) );
  AOI222_X2 U1380 ( .A1(n3138), .A2(n406), .B1(n325), .B2(n403), .C1(n380), 
        .C2(n400), .ZN(n2394) );
  XOR2_X2 U1381 ( .A(n2361), .B(n280), .Z(n1879) );
  OAI21_X4 U1382 ( .B1(n2837), .B2(n354), .A(n2395), .ZN(n2361) );
  AOI222_X2 U1383 ( .A1(n3138), .A2(n403), .B1(n325), .B2(n400), .C1(n380), 
        .C2(n397), .ZN(n2395) );
  XOR2_X2 U1384 ( .A(n2362), .B(n280), .Z(n1880) );
  OAI21_X4 U1385 ( .B1(n2838), .B2(n354), .A(n2396), .ZN(n2362) );
  AOI222_X2 U1386 ( .A1(n3139), .A2(n400), .B1(n325), .B2(n397), .C1(n380), 
        .C2(n393), .ZN(n2396) );
  XOR2_X2 U1387 ( .A(n2363), .B(n280), .Z(n1881) );
  OAI21_X4 U1388 ( .B1(n2839), .B2(n354), .A(n2397), .ZN(n2363) );
  AOI222_X2 U1389 ( .A1(n3138), .A2(n397), .B1(n325), .B2(n393), .C1(n380), 
        .C2(n390), .ZN(n2397) );
  XOR2_X2 U1390 ( .A(n2364), .B(n280), .Z(n1882) );
  OAI21_X4 U1391 ( .B1(n2840), .B2(n354), .A(n2398), .ZN(n2364) );
  XOR2_X2 U1393 ( .A(n2365), .B(n280), .Z(n1883) );
  OAI21_X4 U1394 ( .B1(n2841), .B2(n354), .A(n2399), .ZN(n2365) );
  AND2_X4 U1396 ( .A1(n3138), .A2(n390), .ZN(n1388) );
  XOR2_X2 U1398 ( .A(n2400), .B(n277), .Z(n1885) );
  OAI21_X4 U1399 ( .B1(n2808), .B2(n3130), .A(n2434), .ZN(n2400) );
  NAND2_X4 U1400 ( .A1(n378), .A2(n484), .ZN(n2434) );
  XOR2_X2 U1401 ( .A(n2401), .B(n277), .Z(n1886) );
  OAI21_X4 U1402 ( .B1(n2809), .B2(n3130), .A(n2435), .ZN(n2401) );
  AOI21_X4 U1403 ( .B1(n378), .B2(n481), .A(n1389), .ZN(n2435) );
  AND2_X4 U1404 ( .A1(n323), .A2(n484), .ZN(n1389) );
  XOR2_X2 U1405 ( .A(n2402), .B(n277), .Z(n1887) );
  OAI21_X4 U1406 ( .B1(n2810), .B2(n351), .A(n2436), .ZN(n2402) );
  AOI222_X2 U1407 ( .A1(n3142), .A2(n484), .B1(n323), .B2(n481), .C1(n378), 
        .C2(n478), .ZN(n2436) );
  XOR2_X2 U1408 ( .A(n2403), .B(n277), .Z(n1888) );
  OAI21_X4 U1409 ( .B1(n2811), .B2(n351), .A(n2437), .ZN(n2403) );
  AOI222_X2 U1410 ( .A1(n3141), .A2(n481), .B1(n323), .B2(n478), .C1(n378), 
        .C2(n475), .ZN(n2437) );
  XOR2_X2 U1411 ( .A(n2404), .B(n277), .Z(n1889) );
  OAI21_X4 U1412 ( .B1(n2812), .B2(n351), .A(n2438), .ZN(n2404) );
  AOI222_X2 U1413 ( .A1(n3142), .A2(n478), .B1(n323), .B2(n475), .C1(n378), 
        .C2(n472), .ZN(n2438) );
  XOR2_X2 U1414 ( .A(n2405), .B(n277), .Z(n1890) );
  OAI21_X4 U1415 ( .B1(n2813), .B2(n351), .A(n2439), .ZN(n2405) );
  AOI222_X2 U1416 ( .A1(n3141), .A2(n475), .B1(n323), .B2(n472), .C1(n378), 
        .C2(n469), .ZN(n2439) );
  XOR2_X2 U1417 ( .A(n2406), .B(n277), .Z(n1891) );
  OAI21_X4 U1418 ( .B1(n2814), .B2(n351), .A(n2440), .ZN(n2406) );
  AOI222_X2 U1419 ( .A1(n3142), .A2(n472), .B1(n323), .B2(n469), .C1(n378), 
        .C2(n466), .ZN(n2440) );
  XOR2_X2 U1420 ( .A(n2407), .B(n277), .Z(n1892) );
  OAI21_X4 U1421 ( .B1(n2815), .B2(n351), .A(n2441), .ZN(n2407) );
  AOI222_X2 U1422 ( .A1(n3141), .A2(n469), .B1(n323), .B2(n466), .C1(n378), 
        .C2(n463), .ZN(n2441) );
  XOR2_X2 U1423 ( .A(n2408), .B(n277), .Z(n1893) );
  OAI21_X4 U1424 ( .B1(n2816), .B2(n351), .A(n2442), .ZN(n2408) );
  AOI222_X2 U1425 ( .A1(n3142), .A2(n466), .B1(n323), .B2(n463), .C1(n378), 
        .C2(n460), .ZN(n2442) );
  XOR2_X2 U1426 ( .A(n2409), .B(n277), .Z(n1894) );
  OAI21_X4 U1427 ( .B1(n2817), .B2(n351), .A(n2443), .ZN(n2409) );
  AOI222_X2 U1428 ( .A1(n3141), .A2(n463), .B1(n323), .B2(n460), .C1(n378), 
        .C2(n457), .ZN(n2443) );
  XOR2_X2 U1429 ( .A(n2410), .B(n277), .Z(n1895) );
  OAI21_X4 U1430 ( .B1(n2818), .B2(n351), .A(n2444), .ZN(n2410) );
  AOI222_X2 U1431 ( .A1(n3142), .A2(n460), .B1(n323), .B2(n457), .C1(n378), 
        .C2(n454), .ZN(n2444) );
  XOR2_X2 U1432 ( .A(n2411), .B(n277), .Z(n1896) );
  OAI21_X4 U1433 ( .B1(n2819), .B2(n351), .A(n2445), .ZN(n2411) );
  AOI222_X2 U1434 ( .A1(n3141), .A2(n457), .B1(n323), .B2(n454), .C1(n378), 
        .C2(n451), .ZN(n2445) );
  XOR2_X2 U1435 ( .A(n2412), .B(n277), .Z(n1897) );
  OAI21_X4 U1436 ( .B1(n2820), .B2(n351), .A(n2446), .ZN(n2412) );
  AOI222_X2 U1437 ( .A1(n3141), .A2(n454), .B1(n323), .B2(n451), .C1(n378), 
        .C2(n448), .ZN(n2446) );
  XOR2_X2 U1438 ( .A(n2413), .B(n277), .Z(n1898) );
  OAI21_X4 U1439 ( .B1(n2821), .B2(n351), .A(n2447), .ZN(n2413) );
  AOI222_X2 U1440 ( .A1(n3142), .A2(n451), .B1(n323), .B2(n448), .C1(n378), 
        .C2(n445), .ZN(n2447) );
  XOR2_X2 U1441 ( .A(n2414), .B(n277), .Z(n1899) );
  OAI21_X4 U1442 ( .B1(n2822), .B2(n351), .A(n2448), .ZN(n2414) );
  AOI222_X2 U1443 ( .A1(n3142), .A2(n448), .B1(n323), .B2(n445), .C1(n378), 
        .C2(n442), .ZN(n2448) );
  XOR2_X2 U1444 ( .A(n2415), .B(n277), .Z(n1900) );
  OAI21_X4 U1445 ( .B1(n2823), .B2(n351), .A(n2449), .ZN(n2415) );
  AOI222_X2 U1446 ( .A1(n3142), .A2(n445), .B1(n323), .B2(n442), .C1(n378), 
        .C2(n439), .ZN(n2449) );
  XOR2_X2 U1447 ( .A(n2416), .B(n277), .Z(n1901) );
  OAI21_X4 U1448 ( .B1(n2824), .B2(n351), .A(n2450), .ZN(n2416) );
  AOI222_X2 U1449 ( .A1(n3141), .A2(n442), .B1(n323), .B2(n439), .C1(n378), 
        .C2(n436), .ZN(n2450) );
  XOR2_X2 U1450 ( .A(n2417), .B(n277), .Z(n1902) );
  OAI21_X4 U1451 ( .B1(n2825), .B2(n351), .A(n2451), .ZN(n2417) );
  AOI222_X2 U1452 ( .A1(n3142), .A2(n439), .B1(n323), .B2(n436), .C1(n378), 
        .C2(n433), .ZN(n2451) );
  XOR2_X2 U1453 ( .A(n2418), .B(n277), .Z(n1903) );
  OAI21_X4 U1454 ( .B1(n2826), .B2(n351), .A(n2452), .ZN(n2418) );
  AOI222_X2 U1455 ( .A1(n3141), .A2(n436), .B1(n323), .B2(n433), .C1(n378), 
        .C2(n430), .ZN(n2452) );
  XOR2_X2 U1456 ( .A(n2419), .B(n277), .Z(n1904) );
  OAI21_X4 U1457 ( .B1(n2827), .B2(n351), .A(n2453), .ZN(n2419) );
  AOI222_X2 U1458 ( .A1(n3141), .A2(n433), .B1(n323), .B2(n430), .C1(n378), 
        .C2(n427), .ZN(n2453) );
  XOR2_X2 U1459 ( .A(n2420), .B(n277), .Z(n1905) );
  OAI21_X4 U1460 ( .B1(n2828), .B2(n351), .A(n2454), .ZN(n2420) );
  AOI222_X2 U1461 ( .A1(n3142), .A2(n430), .B1(n323), .B2(n427), .C1(n378), 
        .C2(n424), .ZN(n2454) );
  XOR2_X2 U1462 ( .A(n2421), .B(n277), .Z(n1906) );
  OAI21_X4 U1463 ( .B1(n2829), .B2(n351), .A(n2455), .ZN(n2421) );
  AOI222_X2 U1464 ( .A1(n3141), .A2(n427), .B1(n323), .B2(n424), .C1(n378), 
        .C2(n421), .ZN(n2455) );
  XOR2_X2 U1465 ( .A(n2422), .B(n277), .Z(n1907) );
  OAI21_X4 U1466 ( .B1(n2830), .B2(n351), .A(n2456), .ZN(n2422) );
  AOI222_X2 U1467 ( .A1(n3141), .A2(n424), .B1(n323), .B2(n421), .C1(n378), 
        .C2(n418), .ZN(n2456) );
  XOR2_X2 U1468 ( .A(n2423), .B(n277), .Z(n1908) );
  OAI21_X4 U1469 ( .B1(n2831), .B2(n351), .A(n2457), .ZN(n2423) );
  AOI222_X2 U1470 ( .A1(n3142), .A2(n421), .B1(n323), .B2(n418), .C1(n378), 
        .C2(n415), .ZN(n2457) );
  XOR2_X2 U1471 ( .A(n2424), .B(n277), .Z(n1909) );
  OAI21_X4 U1472 ( .B1(n2832), .B2(n351), .A(n2458), .ZN(n2424) );
  AOI222_X2 U1473 ( .A1(n3142), .A2(n418), .B1(n323), .B2(n415), .C1(n378), 
        .C2(n412), .ZN(n2458) );
  XOR2_X2 U1474 ( .A(n2425), .B(n277), .Z(n1910) );
  OAI21_X4 U1475 ( .B1(n2833), .B2(n351), .A(n2459), .ZN(n2425) );
  AOI222_X2 U1476 ( .A1(n3141), .A2(n415), .B1(n323), .B2(n412), .C1(n378), 
        .C2(n409), .ZN(n2459) );
  XOR2_X2 U1477 ( .A(n2426), .B(n277), .Z(n1911) );
  OAI21_X4 U1478 ( .B1(n2834), .B2(n351), .A(n2460), .ZN(n2426) );
  AOI222_X2 U1479 ( .A1(n3142), .A2(n412), .B1(n323), .B2(n409), .C1(n378), 
        .C2(n406), .ZN(n2460) );
  XOR2_X2 U1480 ( .A(n2427), .B(n277), .Z(n1912) );
  OAI21_X4 U1481 ( .B1(n2835), .B2(n351), .A(n2461), .ZN(n2427) );
  AOI222_X2 U1482 ( .A1(n3141), .A2(n409), .B1(n323), .B2(n406), .C1(n378), 
        .C2(n403), .ZN(n2461) );
  XOR2_X2 U1483 ( .A(n2428), .B(n277), .Z(n1913) );
  OAI21_X4 U1484 ( .B1(n2836), .B2(n351), .A(n2462), .ZN(n2428) );
  AOI222_X2 U1485 ( .A1(n3142), .A2(n406), .B1(n323), .B2(n403), .C1(n378), 
        .C2(n400), .ZN(n2462) );
  XOR2_X2 U1486 ( .A(n2429), .B(n277), .Z(n1914) );
  OAI21_X4 U1487 ( .B1(n2837), .B2(n351), .A(n2463), .ZN(n2429) );
  AOI222_X2 U1488 ( .A1(n3141), .A2(n403), .B1(n323), .B2(n400), .C1(n378), 
        .C2(n397), .ZN(n2463) );
  XOR2_X2 U1489 ( .A(n2430), .B(n277), .Z(n1915) );
  OAI21_X4 U1490 ( .B1(n2838), .B2(n351), .A(n2464), .ZN(n2430) );
  AOI222_X2 U1491 ( .A1(n3142), .A2(n400), .B1(n323), .B2(n397), .C1(n378), 
        .C2(n393), .ZN(n2464) );
  XOR2_X2 U1492 ( .A(n2431), .B(n277), .Z(n1916) );
  OAI21_X4 U1493 ( .B1(n2839), .B2(n351), .A(n2465), .ZN(n2431) );
  AOI222_X2 U1494 ( .A1(n3141), .A2(n397), .B1(n323), .B2(n393), .C1(n378), 
        .C2(n390), .ZN(n2465) );
  XOR2_X2 U1495 ( .A(n2432), .B(n277), .Z(n1917) );
  OAI21_X4 U1496 ( .B1(n2840), .B2(n351), .A(n2466), .ZN(n2432) );
  XOR2_X2 U1498 ( .A(n2433), .B(n277), .Z(n1918) );
  OAI21_X4 U1499 ( .B1(n2841), .B2(n351), .A(n2467), .ZN(n2433) );
  AND2_X4 U1501 ( .A1(n3141), .A2(n390), .ZN(n1391) );
  XOR2_X2 U1503 ( .A(n2468), .B(n274), .Z(n1920) );
  OAI21_X4 U1504 ( .B1(n2808), .B2(n3131), .A(n2502), .ZN(n2468) );
  NAND2_X4 U1505 ( .A1(n376), .A2(n484), .ZN(n2502) );
  XOR2_X2 U1506 ( .A(n2469), .B(n274), .Z(n1921) );
  OAI21_X4 U1507 ( .B1(n2809), .B2(n3131), .A(n2503), .ZN(n2469) );
  AOI21_X4 U1508 ( .B1(n376), .B2(n481), .A(n1392), .ZN(n2503) );
  AND2_X4 U1509 ( .A1(n321), .A2(n484), .ZN(n1392) );
  XOR2_X2 U1510 ( .A(n2470), .B(n274), .Z(n1922) );
  OAI21_X4 U1511 ( .B1(n2810), .B2(n348), .A(n2504), .ZN(n2470) );
  AOI222_X2 U1512 ( .A1(n3185), .A2(n484), .B1(n321), .B2(n481), .C1(n376), 
        .C2(n478), .ZN(n2504) );
  XOR2_X2 U1513 ( .A(n2471), .B(n274), .Z(n1923) );
  OAI21_X4 U1514 ( .B1(n2811), .B2(n348), .A(n2505), .ZN(n2471) );
  AOI222_X2 U1515 ( .A1(n3185), .A2(n481), .B1(n321), .B2(n478), .C1(n376), 
        .C2(n475), .ZN(n2505) );
  XOR2_X2 U1516 ( .A(n2472), .B(n274), .Z(n1924) );
  OAI21_X4 U1517 ( .B1(n2812), .B2(n348), .A(n2506), .ZN(n2472) );
  AOI222_X2 U1518 ( .A1(n3185), .A2(n478), .B1(n321), .B2(n475), .C1(n376), 
        .C2(n472), .ZN(n2506) );
  XOR2_X2 U1519 ( .A(n2473), .B(n274), .Z(n1925) );
  OAI21_X4 U1520 ( .B1(n2813), .B2(n348), .A(n2507), .ZN(n2473) );
  AOI222_X2 U1521 ( .A1(n3185), .A2(n475), .B1(n321), .B2(n472), .C1(n376), 
        .C2(n469), .ZN(n2507) );
  XOR2_X2 U1522 ( .A(n2474), .B(n274), .Z(n1926) );
  OAI21_X4 U1523 ( .B1(n2814), .B2(n348), .A(n2508), .ZN(n2474) );
  AOI222_X2 U1524 ( .A1(n3185), .A2(n472), .B1(n321), .B2(n469), .C1(n376), 
        .C2(n466), .ZN(n2508) );
  XOR2_X2 U1525 ( .A(n2475), .B(n274), .Z(n1927) );
  OAI21_X4 U1526 ( .B1(n2815), .B2(n348), .A(n2509), .ZN(n2475) );
  AOI222_X2 U1527 ( .A1(n3185), .A2(n469), .B1(n321), .B2(n466), .C1(n376), 
        .C2(n463), .ZN(n2509) );
  XOR2_X2 U1528 ( .A(n2476), .B(n274), .Z(n1928) );
  OAI21_X4 U1529 ( .B1(n2816), .B2(n348), .A(n2510), .ZN(n2476) );
  AOI222_X2 U1530 ( .A1(n3185), .A2(n466), .B1(n321), .B2(n463), .C1(n376), 
        .C2(n460), .ZN(n2510) );
  XOR2_X2 U1531 ( .A(n2477), .B(n274), .Z(n1929) );
  OAI21_X4 U1532 ( .B1(n2817), .B2(n348), .A(n2511), .ZN(n2477) );
  AOI222_X2 U1533 ( .A1(n3185), .A2(n463), .B1(n321), .B2(n460), .C1(n376), 
        .C2(n457), .ZN(n2511) );
  XOR2_X2 U1534 ( .A(n2478), .B(n274), .Z(n1930) );
  OAI21_X4 U1535 ( .B1(n2818), .B2(n348), .A(n2512), .ZN(n2478) );
  AOI222_X2 U1536 ( .A1(n3185), .A2(n460), .B1(n321), .B2(n457), .C1(n376), 
        .C2(n454), .ZN(n2512) );
  XOR2_X2 U1537 ( .A(n2479), .B(n274), .Z(n1931) );
  OAI21_X4 U1538 ( .B1(n2819), .B2(n348), .A(n2513), .ZN(n2479) );
  AOI222_X2 U1539 ( .A1(n3185), .A2(n457), .B1(n321), .B2(n454), .C1(n376), 
        .C2(n451), .ZN(n2513) );
  XOR2_X2 U1540 ( .A(n2480), .B(n274), .Z(n1932) );
  OAI21_X4 U1541 ( .B1(n2820), .B2(n348), .A(n2514), .ZN(n2480) );
  AOI222_X2 U1542 ( .A1(n3185), .A2(n454), .B1(n321), .B2(n451), .C1(n376), 
        .C2(n448), .ZN(n2514) );
  XOR2_X2 U1543 ( .A(n2481), .B(n274), .Z(n1933) );
  OAI21_X4 U1544 ( .B1(n2821), .B2(n348), .A(n2515), .ZN(n2481) );
  AOI222_X2 U1545 ( .A1(n3185), .A2(n451), .B1(n321), .B2(n448), .C1(n376), 
        .C2(n445), .ZN(n2515) );
  XOR2_X2 U1546 ( .A(n2482), .B(n274), .Z(n1934) );
  OAI21_X4 U1547 ( .B1(n2822), .B2(n348), .A(n2516), .ZN(n2482) );
  AOI222_X2 U1548 ( .A1(n3185), .A2(n448), .B1(n321), .B2(n445), .C1(n376), 
        .C2(n442), .ZN(n2516) );
  XOR2_X2 U1549 ( .A(n2483), .B(n274), .Z(n1935) );
  OAI21_X4 U1550 ( .B1(n2823), .B2(n348), .A(n2517), .ZN(n2483) );
  AOI222_X2 U1551 ( .A1(n3185), .A2(n445), .B1(n321), .B2(n442), .C1(n376), 
        .C2(n439), .ZN(n2517) );
  XOR2_X2 U1552 ( .A(n2484), .B(n274), .Z(n1936) );
  OAI21_X4 U1553 ( .B1(n2824), .B2(n348), .A(n2518), .ZN(n2484) );
  AOI222_X2 U1554 ( .A1(n3185), .A2(n442), .B1(n321), .B2(n439), .C1(n376), 
        .C2(n436), .ZN(n2518) );
  XOR2_X2 U1555 ( .A(n2485), .B(n274), .Z(n1937) );
  OAI21_X4 U1556 ( .B1(n2825), .B2(n348), .A(n2519), .ZN(n2485) );
  AOI222_X2 U1557 ( .A1(n3185), .A2(n439), .B1(n321), .B2(n436), .C1(n376), 
        .C2(n433), .ZN(n2519) );
  XOR2_X2 U1558 ( .A(n2486), .B(n274), .Z(n1938) );
  OAI21_X4 U1559 ( .B1(n2826), .B2(n348), .A(n2520), .ZN(n2486) );
  AOI222_X2 U1560 ( .A1(n3185), .A2(n436), .B1(n321), .B2(n433), .C1(n376), 
        .C2(n430), .ZN(n2520) );
  XOR2_X2 U1561 ( .A(n2487), .B(n274), .Z(n1939) );
  OAI21_X4 U1562 ( .B1(n2827), .B2(n348), .A(n2521), .ZN(n2487) );
  AOI222_X2 U1563 ( .A1(n3185), .A2(n433), .B1(n321), .B2(n430), .C1(n376), 
        .C2(n427), .ZN(n2521) );
  XOR2_X2 U1564 ( .A(n2488), .B(n274), .Z(n1940) );
  OAI21_X4 U1565 ( .B1(n2828), .B2(n348), .A(n2522), .ZN(n2488) );
  AOI222_X2 U1566 ( .A1(n3185), .A2(n430), .B1(n321), .B2(n427), .C1(n376), 
        .C2(n424), .ZN(n2522) );
  XOR2_X2 U1567 ( .A(n2489), .B(n274), .Z(n1941) );
  OAI21_X4 U1568 ( .B1(n2829), .B2(n348), .A(n2523), .ZN(n2489) );
  AOI222_X2 U1569 ( .A1(n3185), .A2(n427), .B1(n321), .B2(n424), .C1(n376), 
        .C2(n421), .ZN(n2523) );
  XOR2_X2 U1570 ( .A(n2490), .B(n274), .Z(n1942) );
  OAI21_X4 U1571 ( .B1(n2830), .B2(n348), .A(n2524), .ZN(n2490) );
  AOI222_X2 U1572 ( .A1(n3185), .A2(n424), .B1(n321), .B2(n421), .C1(n376), 
        .C2(n418), .ZN(n2524) );
  XOR2_X2 U1573 ( .A(n2491), .B(n274), .Z(n1943) );
  OAI21_X4 U1574 ( .B1(n2831), .B2(n348), .A(n2525), .ZN(n2491) );
  AOI222_X2 U1575 ( .A1(n3185), .A2(n421), .B1(n321), .B2(n418), .C1(n376), 
        .C2(n415), .ZN(n2525) );
  XOR2_X2 U1576 ( .A(n2492), .B(n274), .Z(n1944) );
  OAI21_X4 U1577 ( .B1(n2832), .B2(n348), .A(n2526), .ZN(n2492) );
  AOI222_X2 U1578 ( .A1(n3185), .A2(n418), .B1(n321), .B2(n415), .C1(n376), 
        .C2(n412), .ZN(n2526) );
  XOR2_X2 U1579 ( .A(n2493), .B(n274), .Z(n1945) );
  OAI21_X4 U1580 ( .B1(n2833), .B2(n348), .A(n2527), .ZN(n2493) );
  AOI222_X2 U1581 ( .A1(n3185), .A2(n415), .B1(n321), .B2(n412), .C1(n376), 
        .C2(n409), .ZN(n2527) );
  XOR2_X2 U1582 ( .A(n2494), .B(n274), .Z(n1946) );
  OAI21_X4 U1583 ( .B1(n2834), .B2(n348), .A(n2528), .ZN(n2494) );
  AOI222_X2 U1584 ( .A1(n3185), .A2(n412), .B1(n321), .B2(n409), .C1(n376), 
        .C2(n406), .ZN(n2528) );
  XOR2_X2 U1585 ( .A(n2495), .B(n274), .Z(n1947) );
  OAI21_X4 U1586 ( .B1(n2835), .B2(n348), .A(n2529), .ZN(n2495) );
  AOI222_X2 U1587 ( .A1(n3185), .A2(n409), .B1(n321), .B2(n406), .C1(n376), 
        .C2(n403), .ZN(n2529) );
  XOR2_X2 U1588 ( .A(n2496), .B(n274), .Z(n1948) );
  OAI21_X4 U1589 ( .B1(n2836), .B2(n348), .A(n2530), .ZN(n2496) );
  AOI222_X2 U1590 ( .A1(n3185), .A2(n406), .B1(n321), .B2(n403), .C1(n376), 
        .C2(n400), .ZN(n2530) );
  XOR2_X2 U1591 ( .A(n2497), .B(n274), .Z(n1949) );
  OAI21_X4 U1592 ( .B1(n2837), .B2(n348), .A(n2531), .ZN(n2497) );
  AOI222_X2 U1593 ( .A1(n3185), .A2(n403), .B1(n321), .B2(n400), .C1(n376), 
        .C2(n397), .ZN(n2531) );
  XOR2_X2 U1594 ( .A(n2498), .B(n274), .Z(n1950) );
  OAI21_X4 U1595 ( .B1(n2838), .B2(n348), .A(n2532), .ZN(n2498) );
  AOI222_X2 U1596 ( .A1(n3185), .A2(n400), .B1(n321), .B2(n397), .C1(n376), 
        .C2(n393), .ZN(n2532) );
  XOR2_X2 U1597 ( .A(n2499), .B(n274), .Z(n1951) );
  OAI21_X4 U1598 ( .B1(n2839), .B2(n348), .A(n2533), .ZN(n2499) );
  AOI222_X2 U1599 ( .A1(n3185), .A2(n397), .B1(n321), .B2(n393), .C1(n376), 
        .C2(n390), .ZN(n2533) );
  XOR2_X2 U1600 ( .A(n2500), .B(n274), .Z(n1952) );
  OAI21_X4 U1601 ( .B1(n2840), .B2(n348), .A(n2534), .ZN(n2500) );
  XOR2_X2 U1603 ( .A(n2501), .B(n274), .Z(n1953) );
  OAI21_X4 U1604 ( .B1(n2841), .B2(n348), .A(n2535), .ZN(n2501) );
  AND2_X4 U1606 ( .A1(n3185), .A2(n390), .ZN(n1394) );
  XOR2_X2 U1608 ( .A(n2536), .B(n271), .Z(n1955) );
  OAI21_X4 U1609 ( .B1(n2808), .B2(n3132), .A(n2570), .ZN(n2536) );
  NAND2_X4 U1610 ( .A1(n374), .A2(n484), .ZN(n2570) );
  XOR2_X2 U1611 ( .A(n2537), .B(n271), .Z(n1956) );
  OAI21_X4 U1612 ( .B1(n2809), .B2(n3132), .A(n2571), .ZN(n2537) );
  AOI21_X4 U1613 ( .B1(n374), .B2(n481), .A(n1395), .ZN(n2571) );
  AND2_X4 U1614 ( .A1(n319), .A2(n484), .ZN(n1395) );
  XOR2_X2 U1615 ( .A(n2538), .B(n271), .Z(n1957) );
  OAI21_X4 U1616 ( .B1(n2810), .B2(n345), .A(n2572), .ZN(n2538) );
  AOI222_X2 U1617 ( .A1(n297), .A2(n484), .B1(n319), .B2(n481), .C1(n374), 
        .C2(n478), .ZN(n2572) );
  XOR2_X2 U1618 ( .A(n2539), .B(n271), .Z(n1958) );
  OAI21_X4 U1619 ( .B1(n2811), .B2(n345), .A(n2573), .ZN(n2539) );
  AOI222_X2 U1620 ( .A1(n297), .A2(n481), .B1(n319), .B2(n478), .C1(n374), 
        .C2(n475), .ZN(n2573) );
  XOR2_X2 U1621 ( .A(n2540), .B(n271), .Z(n1959) );
  OAI21_X4 U1622 ( .B1(n2812), .B2(n345), .A(n2574), .ZN(n2540) );
  AOI222_X2 U1623 ( .A1(n297), .A2(n478), .B1(n319), .B2(n475), .C1(n374), 
        .C2(n472), .ZN(n2574) );
  XOR2_X2 U1624 ( .A(n2541), .B(n271), .Z(n1960) );
  OAI21_X4 U1625 ( .B1(n2813), .B2(n345), .A(n2575), .ZN(n2541) );
  AOI222_X2 U1626 ( .A1(n297), .A2(n475), .B1(n319), .B2(n472), .C1(n374), 
        .C2(n469), .ZN(n2575) );
  XOR2_X2 U1627 ( .A(n2542), .B(n271), .Z(n1961) );
  OAI21_X4 U1628 ( .B1(n2814), .B2(n345), .A(n2576), .ZN(n2542) );
  AOI222_X2 U1629 ( .A1(n297), .A2(n472), .B1(n319), .B2(n469), .C1(n374), 
        .C2(n466), .ZN(n2576) );
  XOR2_X2 U1630 ( .A(n2543), .B(n271), .Z(n1962) );
  OAI21_X4 U1631 ( .B1(n2815), .B2(n345), .A(n2577), .ZN(n2543) );
  AOI222_X2 U1632 ( .A1(n297), .A2(n469), .B1(n319), .B2(n466), .C1(n374), 
        .C2(n463), .ZN(n2577) );
  XOR2_X2 U1633 ( .A(n2544), .B(n271), .Z(n1963) );
  OAI21_X4 U1634 ( .B1(n2816), .B2(n345), .A(n2578), .ZN(n2544) );
  AOI222_X2 U1635 ( .A1(n297), .A2(n466), .B1(n319), .B2(n463), .C1(n374), 
        .C2(n460), .ZN(n2578) );
  XOR2_X2 U1636 ( .A(n2545), .B(n271), .Z(n1964) );
  OAI21_X4 U1637 ( .B1(n2817), .B2(n345), .A(n2579), .ZN(n2545) );
  AOI222_X2 U1638 ( .A1(n297), .A2(n463), .B1(n319), .B2(n460), .C1(n374), 
        .C2(n457), .ZN(n2579) );
  XOR2_X2 U1639 ( .A(n2546), .B(n271), .Z(n1965) );
  OAI21_X4 U1640 ( .B1(n2818), .B2(n345), .A(n2580), .ZN(n2546) );
  AOI222_X2 U1641 ( .A1(n297), .A2(n460), .B1(n319), .B2(n457), .C1(n374), 
        .C2(n454), .ZN(n2580) );
  XOR2_X2 U1642 ( .A(n2547), .B(n271), .Z(n1966) );
  OAI21_X4 U1643 ( .B1(n2819), .B2(n345), .A(n2581), .ZN(n2547) );
  AOI222_X2 U1644 ( .A1(n297), .A2(n457), .B1(n319), .B2(n454), .C1(n374), 
        .C2(n451), .ZN(n2581) );
  XOR2_X2 U1645 ( .A(n2548), .B(n271), .Z(n1967) );
  OAI21_X4 U1646 ( .B1(n2820), .B2(n345), .A(n2582), .ZN(n2548) );
  AOI222_X2 U1647 ( .A1(n297), .A2(n454), .B1(n319), .B2(n451), .C1(n374), 
        .C2(n448), .ZN(n2582) );
  XOR2_X2 U1648 ( .A(n2549), .B(n271), .Z(n1968) );
  OAI21_X4 U1649 ( .B1(n2821), .B2(n345), .A(n2583), .ZN(n2549) );
  AOI222_X2 U1650 ( .A1(n297), .A2(n451), .B1(n319), .B2(n448), .C1(n374), 
        .C2(n445), .ZN(n2583) );
  XOR2_X2 U1651 ( .A(n2550), .B(n271), .Z(n1969) );
  OAI21_X4 U1652 ( .B1(n2822), .B2(n345), .A(n2584), .ZN(n2550) );
  AOI222_X2 U1653 ( .A1(n297), .A2(n448), .B1(n319), .B2(n445), .C1(n374), 
        .C2(n442), .ZN(n2584) );
  XOR2_X2 U1654 ( .A(n2551), .B(n271), .Z(n1970) );
  OAI21_X4 U1655 ( .B1(n2823), .B2(n345), .A(n2585), .ZN(n2551) );
  AOI222_X2 U1656 ( .A1(n297), .A2(n445), .B1(n319), .B2(n442), .C1(n374), 
        .C2(n439), .ZN(n2585) );
  XOR2_X2 U1657 ( .A(n2552), .B(n271), .Z(n1971) );
  OAI21_X4 U1658 ( .B1(n2824), .B2(n345), .A(n2586), .ZN(n2552) );
  AOI222_X2 U1659 ( .A1(n297), .A2(n442), .B1(n319), .B2(n439), .C1(n374), 
        .C2(n436), .ZN(n2586) );
  XOR2_X2 U1660 ( .A(n2553), .B(n271), .Z(n1972) );
  OAI21_X4 U1661 ( .B1(n2825), .B2(n345), .A(n2587), .ZN(n2553) );
  AOI222_X2 U1662 ( .A1(n297), .A2(n439), .B1(n319), .B2(n436), .C1(n374), 
        .C2(n433), .ZN(n2587) );
  XOR2_X2 U1663 ( .A(n2554), .B(n271), .Z(n1973) );
  OAI21_X4 U1664 ( .B1(n2826), .B2(n345), .A(n2588), .ZN(n2554) );
  AOI222_X2 U1665 ( .A1(n297), .A2(n436), .B1(n319), .B2(n433), .C1(n374), 
        .C2(n430), .ZN(n2588) );
  XOR2_X2 U1666 ( .A(n2555), .B(n271), .Z(n1974) );
  OAI21_X4 U1667 ( .B1(n2827), .B2(n345), .A(n2589), .ZN(n2555) );
  AOI222_X2 U1668 ( .A1(n297), .A2(n433), .B1(n319), .B2(n430), .C1(n374), 
        .C2(n427), .ZN(n2589) );
  XOR2_X2 U1669 ( .A(n2556), .B(n271), .Z(n1975) );
  OAI21_X4 U1670 ( .B1(n2828), .B2(n345), .A(n2590), .ZN(n2556) );
  AOI222_X2 U1671 ( .A1(n297), .A2(n430), .B1(n319), .B2(n427), .C1(n374), 
        .C2(n424), .ZN(n2590) );
  XOR2_X2 U1672 ( .A(n2557), .B(n271), .Z(n1976) );
  OAI21_X4 U1673 ( .B1(n2829), .B2(n345), .A(n2591), .ZN(n2557) );
  AOI222_X2 U1674 ( .A1(n297), .A2(n427), .B1(n319), .B2(n424), .C1(n374), 
        .C2(n421), .ZN(n2591) );
  XOR2_X2 U1675 ( .A(n2558), .B(n271), .Z(n1977) );
  OAI21_X4 U1676 ( .B1(n2830), .B2(n345), .A(n2592), .ZN(n2558) );
  AOI222_X2 U1677 ( .A1(n297), .A2(n424), .B1(n319), .B2(n421), .C1(n374), 
        .C2(n418), .ZN(n2592) );
  XOR2_X2 U1678 ( .A(n2559), .B(n271), .Z(n1978) );
  OAI21_X4 U1679 ( .B1(n2831), .B2(n345), .A(n2593), .ZN(n2559) );
  AOI222_X2 U1680 ( .A1(n297), .A2(n421), .B1(n319), .B2(n418), .C1(n374), 
        .C2(n415), .ZN(n2593) );
  XOR2_X2 U1681 ( .A(n2560), .B(n271), .Z(n1979) );
  OAI21_X4 U1682 ( .B1(n2832), .B2(n345), .A(n2594), .ZN(n2560) );
  AOI222_X2 U1683 ( .A1(n297), .A2(n418), .B1(n319), .B2(n415), .C1(n374), 
        .C2(n412), .ZN(n2594) );
  XOR2_X2 U1684 ( .A(n2561), .B(n271), .Z(n1980) );
  OAI21_X4 U1685 ( .B1(n2833), .B2(n345), .A(n2595), .ZN(n2561) );
  AOI222_X2 U1686 ( .A1(n297), .A2(n415), .B1(n319), .B2(n412), .C1(n374), 
        .C2(n409), .ZN(n2595) );
  XOR2_X2 U1687 ( .A(n2562), .B(n271), .Z(n1981) );
  OAI21_X4 U1688 ( .B1(n2834), .B2(n345), .A(n2596), .ZN(n2562) );
  AOI222_X2 U1689 ( .A1(n297), .A2(n412), .B1(n319), .B2(n409), .C1(n374), 
        .C2(n406), .ZN(n2596) );
  XOR2_X2 U1690 ( .A(n2563), .B(n271), .Z(n1982) );
  OAI21_X4 U1691 ( .B1(n2835), .B2(n345), .A(n2597), .ZN(n2563) );
  AOI222_X2 U1692 ( .A1(n297), .A2(n409), .B1(n319), .B2(n406), .C1(n374), 
        .C2(n403), .ZN(n2597) );
  XOR2_X2 U1693 ( .A(n2564), .B(n271), .Z(n1983) );
  OAI21_X4 U1694 ( .B1(n2836), .B2(n345), .A(n2598), .ZN(n2564) );
  AOI222_X2 U1695 ( .A1(n297), .A2(n406), .B1(n319), .B2(n403), .C1(n374), 
        .C2(n400), .ZN(n2598) );
  XOR2_X2 U1696 ( .A(n2565), .B(n271), .Z(n1984) );
  OAI21_X4 U1697 ( .B1(n2837), .B2(n345), .A(n2599), .ZN(n2565) );
  AOI222_X2 U1698 ( .A1(n297), .A2(n403), .B1(n319), .B2(n400), .C1(n374), 
        .C2(n397), .ZN(n2599) );
  XOR2_X2 U1699 ( .A(n2566), .B(n271), .Z(n1985) );
  OAI21_X4 U1700 ( .B1(n2838), .B2(n345), .A(n2600), .ZN(n2566) );
  AOI222_X2 U1701 ( .A1(n297), .A2(n400), .B1(n319), .B2(n397), .C1(n374), 
        .C2(n393), .ZN(n2600) );
  XOR2_X2 U1702 ( .A(n2567), .B(n271), .Z(n1986) );
  OAI21_X4 U1703 ( .B1(n2839), .B2(n345), .A(n2601), .ZN(n2567) );
  AOI222_X2 U1704 ( .A1(n297), .A2(n397), .B1(n319), .B2(n393), .C1(n374), 
        .C2(n390), .ZN(n2601) );
  XOR2_X2 U1705 ( .A(n2568), .B(n271), .Z(n1987) );
  OAI21_X4 U1706 ( .B1(n2840), .B2(n345), .A(n2602), .ZN(n2568) );
  OAI21_X4 U1709 ( .B1(n2841), .B2(n345), .A(n2603), .ZN(n2569) );
  AND2_X4 U1711 ( .A1(n297), .A2(n390), .ZN(n1397) );
  XOR2_X2 U1713 ( .A(n2604), .B(n268), .Z(n1990) );
  OAI21_X4 U1714 ( .B1(n2808), .B2(n342), .A(n2638), .ZN(n2604) );
  NAND2_X4 U1715 ( .A1(n3128), .A2(n484), .ZN(n2638) );
  XOR2_X2 U1716 ( .A(n2605), .B(n268), .Z(n1991) );
  OAI21_X4 U1717 ( .B1(n2809), .B2(n342), .A(n2639), .ZN(n2605) );
  AOI21_X4 U1718 ( .B1(n3127), .B2(n481), .A(n1398), .ZN(n2639) );
  AND2_X4 U1719 ( .A1(n317), .A2(n484), .ZN(n1398) );
  XOR2_X2 U1720 ( .A(n2606), .B(n268), .Z(n1992) );
  OAI21_X4 U1721 ( .B1(n2810), .B2(n342), .A(n2640), .ZN(n2606) );
  AOI222_X2 U1722 ( .A1(n295), .A2(n484), .B1(n317), .B2(n481), .C1(n3128), 
        .C2(n478), .ZN(n2640) );
  XOR2_X2 U1723 ( .A(n2607), .B(n268), .Z(n1993) );
  OAI21_X4 U1724 ( .B1(n2811), .B2(n342), .A(n2641), .ZN(n2607) );
  AOI222_X2 U1725 ( .A1(n295), .A2(n481), .B1(n317), .B2(n478), .C1(n3127), 
        .C2(n475), .ZN(n2641) );
  XOR2_X2 U1726 ( .A(n2608), .B(n268), .Z(n1994) );
  OAI21_X4 U1727 ( .B1(n2812), .B2(n342), .A(n2642), .ZN(n2608) );
  AOI222_X2 U1728 ( .A1(n295), .A2(n478), .B1(n317), .B2(n475), .C1(n3128), 
        .C2(n472), .ZN(n2642) );
  XOR2_X2 U1729 ( .A(n2609), .B(n268), .Z(n1995) );
  OAI21_X4 U1730 ( .B1(n2813), .B2(n342), .A(n2643), .ZN(n2609) );
  AOI222_X2 U1731 ( .A1(n295), .A2(n475), .B1(n317), .B2(n472), .C1(n3128), 
        .C2(n469), .ZN(n2643) );
  XOR2_X2 U1732 ( .A(n2610), .B(n268), .Z(n1996) );
  OAI21_X4 U1733 ( .B1(n2814), .B2(n342), .A(n2644), .ZN(n2610) );
  AOI222_X2 U1734 ( .A1(n295), .A2(n472), .B1(n317), .B2(n469), .C1(n3127), 
        .C2(n466), .ZN(n2644) );
  XOR2_X2 U1735 ( .A(n2611), .B(n268), .Z(n1997) );
  OAI21_X4 U1736 ( .B1(n2815), .B2(n342), .A(n2645), .ZN(n2611) );
  AOI222_X2 U1737 ( .A1(n295), .A2(n469), .B1(n317), .B2(n466), .C1(n3128), 
        .C2(n463), .ZN(n2645) );
  XOR2_X2 U1738 ( .A(n2612), .B(n268), .Z(n1998) );
  OAI21_X4 U1739 ( .B1(n2816), .B2(n342), .A(n2646), .ZN(n2612) );
  AOI222_X2 U1740 ( .A1(n295), .A2(n466), .B1(n317), .B2(n463), .C1(n3127), 
        .C2(n460), .ZN(n2646) );
  XOR2_X2 U1741 ( .A(n2613), .B(n268), .Z(n1999) );
  OAI21_X4 U1742 ( .B1(n2817), .B2(n342), .A(n2647), .ZN(n2613) );
  AOI222_X2 U1743 ( .A1(n295), .A2(n463), .B1(n317), .B2(n460), .C1(n3127), 
        .C2(n457), .ZN(n2647) );
  XOR2_X2 U1744 ( .A(n2614), .B(n268), .Z(n2000) );
  OAI21_X4 U1745 ( .B1(n2818), .B2(n342), .A(n2648), .ZN(n2614) );
  AOI222_X2 U1746 ( .A1(n295), .A2(n460), .B1(n317), .B2(n457), .C1(n3128), 
        .C2(n454), .ZN(n2648) );
  XOR2_X2 U1747 ( .A(n2615), .B(n268), .Z(n2001) );
  OAI21_X4 U1748 ( .B1(n2819), .B2(n342), .A(n2649), .ZN(n2615) );
  AOI222_X2 U1749 ( .A1(n295), .A2(n457), .B1(n317), .B2(n454), .C1(n3127), 
        .C2(n451), .ZN(n2649) );
  XOR2_X2 U1750 ( .A(n2616), .B(n268), .Z(n2002) );
  OAI21_X4 U1751 ( .B1(n2820), .B2(n342), .A(n2650), .ZN(n2616) );
  AOI222_X2 U1752 ( .A1(n295), .A2(n454), .B1(n317), .B2(n451), .C1(n3127), 
        .C2(n448), .ZN(n2650) );
  XOR2_X2 U1753 ( .A(n2617), .B(n268), .Z(n2003) );
  OAI21_X4 U1754 ( .B1(n2821), .B2(n342), .A(n2651), .ZN(n2617) );
  AOI222_X2 U1755 ( .A1(n295), .A2(n451), .B1(n317), .B2(n448), .C1(n3128), 
        .C2(n445), .ZN(n2651) );
  XOR2_X2 U1756 ( .A(n2618), .B(n268), .Z(n2004) );
  OAI21_X4 U1757 ( .B1(n2822), .B2(n342), .A(n2652), .ZN(n2618) );
  AOI222_X2 U1758 ( .A1(n295), .A2(n448), .B1(n317), .B2(n445), .C1(n3128), 
        .C2(n442), .ZN(n2652) );
  XOR2_X2 U1759 ( .A(n2619), .B(n268), .Z(n2005) );
  OAI21_X4 U1760 ( .B1(n2823), .B2(n342), .A(n2653), .ZN(n2619) );
  AOI222_X2 U1761 ( .A1(n295), .A2(n445), .B1(n317), .B2(n442), .C1(n3127), 
        .C2(n439), .ZN(n2653) );
  XOR2_X2 U1762 ( .A(n2620), .B(n268), .Z(n2006) );
  OAI21_X4 U1763 ( .B1(n2824), .B2(n342), .A(n2654), .ZN(n2620) );
  AOI222_X2 U1764 ( .A1(n295), .A2(n442), .B1(n317), .B2(n439), .C1(n3128), 
        .C2(n436), .ZN(n2654) );
  XOR2_X2 U1765 ( .A(n2621), .B(n268), .Z(n2007) );
  OAI21_X4 U1766 ( .B1(n2825), .B2(n342), .A(n2655), .ZN(n2621) );
  AOI222_X2 U1767 ( .A1(n295), .A2(n439), .B1(n317), .B2(n436), .C1(n3127), 
        .C2(n433), .ZN(n2655) );
  XOR2_X2 U1768 ( .A(n2622), .B(n268), .Z(n2008) );
  OAI21_X4 U1769 ( .B1(n2826), .B2(n342), .A(n2656), .ZN(n2622) );
  AOI222_X2 U1770 ( .A1(n295), .A2(n436), .B1(n317), .B2(n433), .C1(n3128), 
        .C2(n430), .ZN(n2656) );
  XOR2_X2 U1771 ( .A(n2623), .B(n268), .Z(n2009) );
  OAI21_X4 U1772 ( .B1(n2827), .B2(n342), .A(n2657), .ZN(n2623) );
  AOI222_X2 U1773 ( .A1(n295), .A2(n433), .B1(n317), .B2(n430), .C1(n3128), 
        .C2(n427), .ZN(n2657) );
  XOR2_X2 U1774 ( .A(n2624), .B(n268), .Z(n2010) );
  OAI21_X4 U1775 ( .B1(n2828), .B2(n342), .A(n2658), .ZN(n2624) );
  AOI222_X2 U1776 ( .A1(n295), .A2(n430), .B1(n317), .B2(n427), .C1(n3127), 
        .C2(n424), .ZN(n2658) );
  XOR2_X2 U1777 ( .A(n2625), .B(n268), .Z(n2011) );
  OAI21_X4 U1778 ( .B1(n2829), .B2(n342), .A(n2659), .ZN(n2625) );
  AOI222_X2 U1779 ( .A1(n295), .A2(n427), .B1(n317), .B2(n424), .C1(n3128), 
        .C2(n421), .ZN(n2659) );
  XOR2_X2 U1780 ( .A(n2626), .B(n268), .Z(n2012) );
  OAI21_X4 U1781 ( .B1(n2830), .B2(n342), .A(n2660), .ZN(n2626) );
  AOI222_X2 U1782 ( .A1(n295), .A2(n424), .B1(n317), .B2(n421), .C1(n3127), 
        .C2(n418), .ZN(n2660) );
  XOR2_X2 U1783 ( .A(n2627), .B(n268), .Z(n2013) );
  OAI21_X4 U1784 ( .B1(n2831), .B2(n342), .A(n2661), .ZN(n2627) );
  AOI222_X2 U1785 ( .A1(n295), .A2(n421), .B1(n317), .B2(n418), .C1(n3128), 
        .C2(n415), .ZN(n2661) );
  XOR2_X2 U1786 ( .A(n2628), .B(n268), .Z(n2014) );
  OAI21_X4 U1787 ( .B1(n2832), .B2(n342), .A(n2662), .ZN(n2628) );
  AOI222_X2 U1788 ( .A1(n295), .A2(n418), .B1(n317), .B2(n415), .C1(n3127), 
        .C2(n412), .ZN(n2662) );
  XOR2_X2 U1789 ( .A(n2629), .B(n268), .Z(n2015) );
  OAI21_X4 U1790 ( .B1(n2833), .B2(n342), .A(n2663), .ZN(n2629) );
  AOI222_X2 U1791 ( .A1(n295), .A2(n415), .B1(n317), .B2(n412), .C1(n3127), 
        .C2(n409), .ZN(n2663) );
  XOR2_X2 U1792 ( .A(n2630), .B(n268), .Z(n2016) );
  OAI21_X4 U1793 ( .B1(n2834), .B2(n342), .A(n2664), .ZN(n2630) );
  AOI222_X2 U1794 ( .A1(n295), .A2(n412), .B1(n317), .B2(n409), .C1(n3127), 
        .C2(n406), .ZN(n2664) );
  XOR2_X2 U1795 ( .A(n2631), .B(n268), .Z(n2017) );
  OAI21_X4 U1796 ( .B1(n2835), .B2(n342), .A(n2665), .ZN(n2631) );
  AOI222_X2 U1797 ( .A1(n295), .A2(n409), .B1(n317), .B2(n406), .C1(n3128), 
        .C2(n403), .ZN(n2665) );
  XOR2_X2 U1798 ( .A(n2632), .B(n268), .Z(n2018) );
  OAI21_X4 U1799 ( .B1(n2836), .B2(n342), .A(n2666), .ZN(n2632) );
  AOI222_X2 U1800 ( .A1(n295), .A2(n406), .B1(n317), .B2(n403), .C1(n3128), 
        .C2(n400), .ZN(n2666) );
  XOR2_X2 U1801 ( .A(n2633), .B(n268), .Z(n2019) );
  OAI21_X4 U1802 ( .B1(n2837), .B2(n342), .A(n2667), .ZN(n2633) );
  AOI222_X2 U1803 ( .A1(n295), .A2(n403), .B1(n317), .B2(n400), .C1(n3127), 
        .C2(n397), .ZN(n2667) );
  XOR2_X2 U1804 ( .A(n2634), .B(n268), .Z(n2020) );
  OAI21_X4 U1805 ( .B1(n2838), .B2(n342), .A(n2668), .ZN(n2634) );
  AOI222_X2 U1806 ( .A1(n295), .A2(n400), .B1(n317), .B2(n397), .C1(n3128), 
        .C2(n393), .ZN(n2668) );
  XOR2_X2 U1807 ( .A(n2635), .B(n268), .Z(n2021) );
  XOR2_X2 U1810 ( .A(n2636), .B(n268), .Z(n2022) );
  AND2_X4 U1816 ( .A1(n295), .A2(n390), .ZN(n1400) );
  XOR2_X2 U1818 ( .A(n2672), .B(n265), .Z(n2025) );
  OAI21_X4 U1819 ( .B1(n2808), .B2(n339), .A(n2706), .ZN(n2672) );
  NAND2_X4 U1820 ( .A1(n370), .A2(n484), .ZN(n2706) );
  XOR2_X2 U1821 ( .A(n2673), .B(n265), .Z(n2026) );
  OAI21_X4 U1822 ( .B1(n2809), .B2(n339), .A(n2707), .ZN(n2673) );
  AOI21_X4 U1823 ( .B1(n370), .B2(n481), .A(n1401), .ZN(n2707) );
  AND2_X4 U1824 ( .A1(n315), .A2(n484), .ZN(n1401) );
  XOR2_X2 U1825 ( .A(n2674), .B(n265), .Z(n2027) );
  OAI21_X4 U1826 ( .B1(n2810), .B2(n339), .A(n2708), .ZN(n2674) );
  AOI222_X2 U1827 ( .A1(n293), .A2(n484), .B1(n315), .B2(n481), .C1(n370), 
        .C2(n478), .ZN(n2708) );
  XOR2_X2 U1828 ( .A(n2675), .B(n265), .Z(n2028) );
  OAI21_X4 U1829 ( .B1(n2811), .B2(n339), .A(n2709), .ZN(n2675) );
  AOI222_X2 U1830 ( .A1(n293), .A2(n481), .B1(n315), .B2(n478), .C1(n370), 
        .C2(n475), .ZN(n2709) );
  XOR2_X2 U1831 ( .A(n2676), .B(n265), .Z(n2029) );
  OAI21_X4 U1832 ( .B1(n2812), .B2(n339), .A(n2710), .ZN(n2676) );
  AOI222_X2 U1833 ( .A1(n293), .A2(n478), .B1(n315), .B2(n475), .C1(n370), 
        .C2(n472), .ZN(n2710) );
  XOR2_X2 U1834 ( .A(n2677), .B(n265), .Z(n2030) );
  OAI21_X4 U1835 ( .B1(n2813), .B2(n339), .A(n2711), .ZN(n2677) );
  AOI222_X2 U1836 ( .A1(n293), .A2(n475), .B1(n315), .B2(n472), .C1(n370), 
        .C2(n469), .ZN(n2711) );
  XOR2_X2 U1837 ( .A(n2678), .B(n265), .Z(n2031) );
  OAI21_X4 U1838 ( .B1(n2814), .B2(n339), .A(n2712), .ZN(n2678) );
  AOI222_X2 U1839 ( .A1(n293), .A2(n472), .B1(n315), .B2(n469), .C1(n370), 
        .C2(n466), .ZN(n2712) );
  XOR2_X2 U1840 ( .A(n2679), .B(n265), .Z(n2032) );
  OAI21_X4 U1841 ( .B1(n2815), .B2(n339), .A(n2713), .ZN(n2679) );
  AOI222_X2 U1842 ( .A1(n293), .A2(n469), .B1(n315), .B2(n466), .C1(n370), 
        .C2(n463), .ZN(n2713) );
  XOR2_X2 U1843 ( .A(n2680), .B(n265), .Z(n2033) );
  OAI21_X4 U1844 ( .B1(n2816), .B2(n339), .A(n2714), .ZN(n2680) );
  AOI222_X2 U1845 ( .A1(n293), .A2(n466), .B1(n315), .B2(n463), .C1(n370), 
        .C2(n460), .ZN(n2714) );
  XOR2_X2 U1846 ( .A(n2681), .B(n265), .Z(n2034) );
  OAI21_X4 U1847 ( .B1(n2817), .B2(n339), .A(n2715), .ZN(n2681) );
  AOI222_X2 U1848 ( .A1(n293), .A2(n463), .B1(n315), .B2(n460), .C1(n370), 
        .C2(n457), .ZN(n2715) );
  XOR2_X2 U1849 ( .A(n2682), .B(n265), .Z(n2035) );
  OAI21_X4 U1850 ( .B1(n2818), .B2(n339), .A(n2716), .ZN(n2682) );
  AOI222_X2 U1851 ( .A1(n293), .A2(n460), .B1(n315), .B2(n457), .C1(n370), 
        .C2(n454), .ZN(n2716) );
  XOR2_X2 U1852 ( .A(n2683), .B(n265), .Z(n2036) );
  OAI21_X4 U1853 ( .B1(n2819), .B2(n339), .A(n2717), .ZN(n2683) );
  AOI222_X2 U1854 ( .A1(n293), .A2(n457), .B1(n315), .B2(n454), .C1(n370), 
        .C2(n451), .ZN(n2717) );
  XOR2_X2 U1855 ( .A(n2684), .B(n265), .Z(n2037) );
  OAI21_X4 U1856 ( .B1(n2820), .B2(n339), .A(n2718), .ZN(n2684) );
  AOI222_X2 U1857 ( .A1(n293), .A2(n454), .B1(n315), .B2(n451), .C1(n370), 
        .C2(n448), .ZN(n2718) );
  XOR2_X2 U1858 ( .A(n2685), .B(n265), .Z(n2038) );
  OAI21_X4 U1859 ( .B1(n2821), .B2(n339), .A(n2719), .ZN(n2685) );
  AOI222_X2 U1860 ( .A1(n293), .A2(n451), .B1(n315), .B2(n448), .C1(n370), 
        .C2(n445), .ZN(n2719) );
  XOR2_X2 U1861 ( .A(n2686), .B(n265), .Z(n2039) );
  OAI21_X4 U1862 ( .B1(n2822), .B2(n339), .A(n2720), .ZN(n2686) );
  AOI222_X2 U1863 ( .A1(n293), .A2(n448), .B1(n315), .B2(n445), .C1(n370), 
        .C2(n442), .ZN(n2720) );
  XOR2_X2 U1864 ( .A(n2687), .B(n265), .Z(n2040) );
  OAI21_X4 U1865 ( .B1(n2823), .B2(n339), .A(n2721), .ZN(n2687) );
  AOI222_X2 U1866 ( .A1(n293), .A2(n445), .B1(n315), .B2(n442), .C1(n370), 
        .C2(n439), .ZN(n2721) );
  XOR2_X2 U1867 ( .A(n2688), .B(n265), .Z(n2041) );
  OAI21_X4 U1868 ( .B1(n2824), .B2(n339), .A(n2722), .ZN(n2688) );
  AOI222_X2 U1869 ( .A1(n293), .A2(n442), .B1(n315), .B2(n439), .C1(n370), 
        .C2(n436), .ZN(n2722) );
  XOR2_X2 U1870 ( .A(n2689), .B(n265), .Z(n2042) );
  OAI21_X4 U1871 ( .B1(n2825), .B2(n339), .A(n2723), .ZN(n2689) );
  AOI222_X2 U1872 ( .A1(n293), .A2(n439), .B1(n315), .B2(n436), .C1(n370), 
        .C2(n433), .ZN(n2723) );
  XOR2_X2 U1873 ( .A(n2690), .B(n265), .Z(n2043) );
  OAI21_X4 U1874 ( .B1(n2826), .B2(n339), .A(n2724), .ZN(n2690) );
  AOI222_X2 U1875 ( .A1(n293), .A2(n436), .B1(n315), .B2(n433), .C1(n370), 
        .C2(n430), .ZN(n2724) );
  XOR2_X2 U1876 ( .A(n2691), .B(n265), .Z(n2044) );
  OAI21_X4 U1877 ( .B1(n2827), .B2(n339), .A(n2725), .ZN(n2691) );
  AOI222_X2 U1878 ( .A1(n293), .A2(n433), .B1(n315), .B2(n430), .C1(n370), 
        .C2(n427), .ZN(n2725) );
  XOR2_X2 U1879 ( .A(n2692), .B(n265), .Z(n2045) );
  OAI21_X4 U1880 ( .B1(n2828), .B2(n339), .A(n2726), .ZN(n2692) );
  AOI222_X2 U1881 ( .A1(n293), .A2(n430), .B1(n315), .B2(n427), .C1(n370), 
        .C2(n424), .ZN(n2726) );
  XOR2_X2 U1882 ( .A(n2693), .B(n265), .Z(n2046) );
  OAI21_X4 U1883 ( .B1(n2829), .B2(n339), .A(n2727), .ZN(n2693) );
  AOI222_X2 U1884 ( .A1(n293), .A2(n427), .B1(n315), .B2(n424), .C1(n370), 
        .C2(n421), .ZN(n2727) );
  XOR2_X2 U1885 ( .A(n2694), .B(n265), .Z(n2047) );
  OAI21_X4 U1886 ( .B1(n2830), .B2(n339), .A(n2728), .ZN(n2694) );
  AOI222_X2 U1887 ( .A1(n293), .A2(n424), .B1(n315), .B2(n421), .C1(n370), 
        .C2(n418), .ZN(n2728) );
  XOR2_X2 U1888 ( .A(n2695), .B(n265), .Z(n2048) );
  OAI21_X4 U1889 ( .B1(n2831), .B2(n339), .A(n2729), .ZN(n2695) );
  AOI222_X2 U1890 ( .A1(n293), .A2(n421), .B1(n315), .B2(n418), .C1(n370), 
        .C2(n415), .ZN(n2729) );
  XOR2_X2 U1891 ( .A(n2696), .B(n265), .Z(n2049) );
  OAI21_X4 U1892 ( .B1(n2832), .B2(n339), .A(n2730), .ZN(n2696) );
  AOI222_X2 U1893 ( .A1(n293), .A2(n418), .B1(n315), .B2(n415), .C1(n370), 
        .C2(n412), .ZN(n2730) );
  XOR2_X2 U1894 ( .A(n2697), .B(n265), .Z(n2050) );
  OAI21_X4 U1895 ( .B1(n2833), .B2(n339), .A(n2731), .ZN(n2697) );
  AOI222_X2 U1896 ( .A1(n293), .A2(n415), .B1(n315), .B2(n412), .C1(n370), 
        .C2(n409), .ZN(n2731) );
  XOR2_X2 U1897 ( .A(n2698), .B(n265), .Z(n2051) );
  OAI21_X4 U1898 ( .B1(n2834), .B2(n339), .A(n2732), .ZN(n2698) );
  AOI222_X2 U1899 ( .A1(n293), .A2(n412), .B1(n315), .B2(n409), .C1(n370), 
        .C2(n406), .ZN(n2732) );
  XOR2_X2 U1900 ( .A(n2699), .B(n265), .Z(n2052) );
  OAI21_X4 U1901 ( .B1(n2835), .B2(n339), .A(n2733), .ZN(n2699) );
  AOI222_X2 U1902 ( .A1(n293), .A2(n409), .B1(n315), .B2(n406), .C1(n370), 
        .C2(n403), .ZN(n2733) );
  XOR2_X2 U1903 ( .A(n2700), .B(n265), .Z(n2053) );
  OAI21_X4 U1904 ( .B1(n2836), .B2(n339), .A(n2734), .ZN(n2700) );
  AOI222_X2 U1905 ( .A1(n293), .A2(n406), .B1(n315), .B2(n403), .C1(n370), 
        .C2(n400), .ZN(n2734) );
  XOR2_X2 U1906 ( .A(n2701), .B(n265), .Z(n2054) );
  OAI21_X4 U1907 ( .B1(n2837), .B2(n339), .A(n2735), .ZN(n2701) );
  AOI222_X2 U1908 ( .A1(n293), .A2(n403), .B1(n315), .B2(n400), .C1(n370), 
        .C2(n397), .ZN(n2735) );
  XOR2_X2 U1909 ( .A(n2702), .B(n265), .Z(n2055) );
  OAI21_X4 U1910 ( .B1(n2838), .B2(n339), .A(n2736), .ZN(n2702) );
  AOI222_X2 U1911 ( .A1(n293), .A2(n400), .B1(n315), .B2(n397), .C1(n370), 
        .C2(n393), .ZN(n2736) );
  XOR2_X2 U1912 ( .A(n2703), .B(n265), .Z(n2056) );
  OAI21_X4 U1913 ( .B1(n2839), .B2(n339), .A(n2737), .ZN(n2703) );
  AOI222_X2 U1914 ( .A1(n293), .A2(n397), .B1(n315), .B2(n393), .C1(n370), 
        .C2(n390), .ZN(n2737) );
  XOR2_X2 U1915 ( .A(n2704), .B(n265), .Z(n2057) );
  OAI21_X4 U1919 ( .B1(n2841), .B2(n339), .A(n2739), .ZN(n2705) );
  AND2_X4 U1921 ( .A1(n293), .A2(n390), .ZN(n1403) );
  XOR2_X2 U1923 ( .A(n2740), .B(n262), .Z(n2060) );
  OAI21_X4 U1924 ( .B1(n2808), .B2(n3133), .A(n2774), .ZN(n2740) );
  NAND2_X4 U1925 ( .A1(n368), .A2(n484), .ZN(n2774) );
  XOR2_X2 U1926 ( .A(n2741), .B(n262), .Z(n2061) );
  OAI21_X4 U1927 ( .B1(n2809), .B2(n3133), .A(n2775), .ZN(n2741) );
  AOI21_X4 U1928 ( .B1(n368), .B2(n481), .A(n1404), .ZN(n2775) );
  AND2_X4 U1929 ( .A1(n313), .A2(n484), .ZN(n1404) );
  XOR2_X2 U1930 ( .A(n2742), .B(n262), .Z(n2062) );
  OAI21_X4 U1931 ( .B1(n2810), .B2(n3133), .A(n2776), .ZN(n2742) );
  AOI222_X2 U1932 ( .A1(n3154), .A2(n484), .B1(n313), .B2(n481), .C1(n368), 
        .C2(n478), .ZN(n2776) );
  XOR2_X2 U1933 ( .A(n2743), .B(n262), .Z(n2063) );
  OAI21_X4 U1934 ( .B1(n2811), .B2(n336), .A(n2777), .ZN(n2743) );
  AOI222_X2 U1935 ( .A1(n3154), .A2(n481), .B1(n313), .B2(n478), .C1(n368), 
        .C2(n475), .ZN(n2777) );
  XOR2_X2 U1936 ( .A(n2744), .B(n262), .Z(n2064) );
  OAI21_X4 U1937 ( .B1(n2812), .B2(n336), .A(n2778), .ZN(n2744) );
  AOI222_X2 U1938 ( .A1(n3153), .A2(n478), .B1(n313), .B2(n475), .C1(n368), 
        .C2(n472), .ZN(n2778) );
  XOR2_X2 U1939 ( .A(n2745), .B(n262), .Z(n2065) );
  OAI21_X4 U1940 ( .B1(n2813), .B2(n336), .A(n2779), .ZN(n2745) );
  AOI222_X2 U1941 ( .A1(n3153), .A2(n475), .B1(n313), .B2(n472), .C1(n368), 
        .C2(n469), .ZN(n2779) );
  XOR2_X2 U1942 ( .A(n2746), .B(n262), .Z(n2066) );
  OAI21_X4 U1943 ( .B1(n2814), .B2(n336), .A(n2780), .ZN(n2746) );
  AOI222_X2 U1944 ( .A1(n3153), .A2(n472), .B1(n313), .B2(n469), .C1(n368), 
        .C2(n466), .ZN(n2780) );
  XOR2_X2 U1945 ( .A(n2747), .B(n262), .Z(n2067) );
  OAI21_X4 U1946 ( .B1(n2815), .B2(n336), .A(n2781), .ZN(n2747) );
  AOI222_X2 U1947 ( .A1(n3154), .A2(n469), .B1(n313), .B2(n466), .C1(n368), 
        .C2(n463), .ZN(n2781) );
  XOR2_X2 U1948 ( .A(n2748), .B(n262), .Z(n2068) );
  OAI21_X4 U1949 ( .B1(n2816), .B2(n336), .A(n2782), .ZN(n2748) );
  AOI222_X2 U1950 ( .A1(n3154), .A2(n466), .B1(n313), .B2(n463), .C1(n368), 
        .C2(n460), .ZN(n2782) );
  XOR2_X2 U1951 ( .A(n2749), .B(n262), .Z(n2069) );
  OAI21_X4 U1952 ( .B1(n2817), .B2(n336), .A(n2783), .ZN(n2749) );
  AOI222_X2 U1953 ( .A1(n3153), .A2(n463), .B1(n313), .B2(n460), .C1(n368), 
        .C2(n457), .ZN(n2783) );
  XOR2_X2 U1954 ( .A(n2750), .B(n262), .Z(n2070) );
  OAI21_X4 U1955 ( .B1(n2818), .B2(n336), .A(n2784), .ZN(n2750) );
  AOI222_X2 U1956 ( .A1(n3154), .A2(n460), .B1(n313), .B2(n457), .C1(n368), 
        .C2(n454), .ZN(n2784) );
  XOR2_X2 U1957 ( .A(n2751), .B(n262), .Z(n2071) );
  OAI21_X4 U1958 ( .B1(n2819), .B2(n336), .A(n2785), .ZN(n2751) );
  AOI222_X2 U1959 ( .A1(n3153), .A2(n457), .B1(n313), .B2(n454), .C1(n368), 
        .C2(n451), .ZN(n2785) );
  XOR2_X2 U1960 ( .A(n2752), .B(n262), .Z(n2072) );
  OAI21_X4 U1961 ( .B1(n2820), .B2(n336), .A(n2786), .ZN(n2752) );
  AOI222_X2 U1962 ( .A1(n3154), .A2(n454), .B1(n313), .B2(n451), .C1(n368), 
        .C2(n448), .ZN(n2786) );
  XOR2_X2 U1963 ( .A(n2753), .B(n262), .Z(n2073) );
  OAI21_X4 U1964 ( .B1(n2821), .B2(n336), .A(n2787), .ZN(n2753) );
  AOI222_X2 U1965 ( .A1(n3153), .A2(n451), .B1(n313), .B2(n448), .C1(n368), 
        .C2(n445), .ZN(n2787) );
  XOR2_X2 U1966 ( .A(n2754), .B(n262), .Z(n2074) );
  OAI21_X4 U1967 ( .B1(n2822), .B2(n336), .A(n2788), .ZN(n2754) );
  AOI222_X2 U1968 ( .A1(n3154), .A2(n448), .B1(n313), .B2(n445), .C1(n368), 
        .C2(n442), .ZN(n2788) );
  XOR2_X2 U1969 ( .A(n2755), .B(n262), .Z(n2075) );
  OAI21_X4 U1970 ( .B1(n2823), .B2(n336), .A(n2789), .ZN(n2755) );
  AOI222_X2 U1971 ( .A1(n3153), .A2(n445), .B1(n313), .B2(n442), .C1(n368), 
        .C2(n439), .ZN(n2789) );
  XOR2_X2 U1972 ( .A(n2756), .B(n262), .Z(n2076) );
  OAI21_X4 U1973 ( .B1(n2824), .B2(n336), .A(n2790), .ZN(n2756) );
  AOI222_X2 U1974 ( .A1(n3154), .A2(n442), .B1(n313), .B2(n439), .C1(n368), 
        .C2(n436), .ZN(n2790) );
  XOR2_X2 U1975 ( .A(n2757), .B(n262), .Z(n2077) );
  OAI21_X4 U1976 ( .B1(n2825), .B2(n336), .A(n2791), .ZN(n2757) );
  AOI222_X2 U1977 ( .A1(n3153), .A2(n439), .B1(n313), .B2(n436), .C1(n368), 
        .C2(n433), .ZN(n2791) );
  XOR2_X2 U1978 ( .A(n2758), .B(n262), .Z(n2078) );
  OAI21_X4 U1979 ( .B1(n2826), .B2(n336), .A(n2792), .ZN(n2758) );
  AOI222_X2 U1980 ( .A1(n3153), .A2(n436), .B1(n313), .B2(n433), .C1(n368), 
        .C2(n430), .ZN(n2792) );
  XOR2_X2 U1981 ( .A(n2759), .B(n262), .Z(n2079) );
  OAI21_X4 U1982 ( .B1(n2827), .B2(n336), .A(n2793), .ZN(n2759) );
  AOI222_X2 U1983 ( .A1(n3154), .A2(n433), .B1(n313), .B2(n430), .C1(n368), 
        .C2(n427), .ZN(n2793) );
  XOR2_X2 U1984 ( .A(n2760), .B(n262), .Z(n2080) );
  OAI21_X4 U1985 ( .B1(n2828), .B2(n336), .A(n2794), .ZN(n2760) );
  AOI222_X2 U1986 ( .A1(n3154), .A2(n430), .B1(n313), .B2(n427), .C1(n368), 
        .C2(n424), .ZN(n2794) );
  XOR2_X2 U1987 ( .A(n2761), .B(n262), .Z(n2081) );
  OAI21_X4 U1988 ( .B1(n2829), .B2(n336), .A(n2795), .ZN(n2761) );
  AOI222_X2 U1989 ( .A1(n3154), .A2(n427), .B1(n313), .B2(n424), .C1(n368), 
        .C2(n421), .ZN(n2795) );
  XOR2_X2 U1990 ( .A(n2762), .B(n262), .Z(n2082) );
  OAI21_X4 U1991 ( .B1(n2830), .B2(n336), .A(n2796), .ZN(n2762) );
  AOI222_X2 U1992 ( .A1(n3154), .A2(n424), .B1(n313), .B2(n421), .C1(n368), 
        .C2(n418), .ZN(n2796) );
  XOR2_X2 U1993 ( .A(n2763), .B(n262), .Z(n2083) );
  OAI21_X4 U1994 ( .B1(n2831), .B2(n336), .A(n2797), .ZN(n2763) );
  AOI222_X2 U1995 ( .A1(n3153), .A2(n421), .B1(n313), .B2(n418), .C1(n368), 
        .C2(n415), .ZN(n2797) );
  XOR2_X2 U1996 ( .A(n2764), .B(n262), .Z(n2084) );
  OAI21_X4 U1997 ( .B1(n2832), .B2(n336), .A(n2798), .ZN(n2764) );
  AOI222_X2 U1998 ( .A1(n3154), .A2(n418), .B1(n313), .B2(n415), .C1(n368), 
        .C2(n412), .ZN(n2798) );
  XOR2_X2 U1999 ( .A(n2765), .B(n262), .Z(n2085) );
  OAI21_X4 U2000 ( .B1(n2833), .B2(n336), .A(n2799), .ZN(n2765) );
  AOI222_X2 U2001 ( .A1(n3153), .A2(n415), .B1(n313), .B2(n412), .C1(n368), 
        .C2(n409), .ZN(n2799) );
  XOR2_X2 U2002 ( .A(n2766), .B(n262), .Z(n2086) );
  OAI21_X4 U2003 ( .B1(n2834), .B2(n336), .A(n2800), .ZN(n2766) );
  AOI222_X2 U2004 ( .A1(n3153), .A2(n412), .B1(n313), .B2(n409), .C1(n368), 
        .C2(n406), .ZN(n2800) );
  XOR2_X2 U2005 ( .A(n2767), .B(n262), .Z(n2087) );
  OAI21_X4 U2006 ( .B1(n2835), .B2(n336), .A(n2801), .ZN(n2767) );
  AOI222_X2 U2007 ( .A1(n3153), .A2(n409), .B1(n313), .B2(n406), .C1(n368), 
        .C2(n403), .ZN(n2801) );
  XOR2_X2 U2008 ( .A(n2768), .B(n262), .Z(n2088) );
  OAI21_X4 U2009 ( .B1(n2836), .B2(n336), .A(n2802), .ZN(n2768) );
  AOI222_X2 U2010 ( .A1(n3153), .A2(n406), .B1(n313), .B2(n403), .C1(n368), 
        .C2(n400), .ZN(n2802) );
  XOR2_X2 U2011 ( .A(n2769), .B(n262), .Z(n2089) );
  OAI21_X4 U2012 ( .B1(n2837), .B2(n336), .A(n2803), .ZN(n2769) );
  AOI222_X2 U2013 ( .A1(n3154), .A2(n403), .B1(n313), .B2(n400), .C1(n368), 
        .C2(n397), .ZN(n2803) );
  XOR2_X2 U2014 ( .A(n2770), .B(n262), .Z(n2090) );
  OAI21_X4 U2015 ( .B1(n2838), .B2(n336), .A(n2804), .ZN(n2770) );
  AOI222_X2 U2016 ( .A1(n3154), .A2(n400), .B1(n313), .B2(n397), .C1(n368), 
        .C2(n393), .ZN(n2804) );
  XOR2_X2 U2017 ( .A(n2771), .B(n262), .Z(n2091) );
  OAI21_X4 U2018 ( .B1(n2839), .B2(n336), .A(n2805), .ZN(n2771) );
  AOI222_X2 U2019 ( .A1(n3153), .A2(n397), .B1(n313), .B2(n393), .C1(n368), 
        .C2(n390), .ZN(n2805) );
  XOR2_X2 U2020 ( .A(n2772), .B(n262), .Z(n678) );
  OAI21_X4 U2021 ( .B1(n2840), .B2(n336), .A(n2806), .ZN(n2772) );
  XOR2_X2 U2023 ( .A(n2773), .B(n262), .Z(n2093) );
  OAI21_X4 U2024 ( .B1(n2841), .B2(n336), .A(n2807), .ZN(n2773) );
  AND2_X4 U2026 ( .A1(n3153), .A2(n390), .ZN(n1406) );
  AND3_X4 U2103 ( .A1(n2908), .A2(n2919), .A3(a[31]), .ZN(n388) );
  AND3_X4 U2107 ( .A1(n2931), .A2(n2909), .A3(n2920), .ZN(n386) );
  AND3_X4 U2112 ( .A1(n2932), .A2(n2910), .A3(n2921), .ZN(n384) );
  AND3_X4 U2117 ( .A1(n2933), .A2(n2911), .A3(n2922), .ZN(n382) );
  AND3_X4 U2122 ( .A1(n2934), .A2(n2912), .A3(n2923), .ZN(n380) );
  AND3_X4 U2127 ( .A1(n2935), .A2(n2913), .A3(n2924), .ZN(n378) );
  AND3_X4 U2132 ( .A1(n2936), .A2(n2914), .A3(n2925), .ZN(n376) );
  XNOR2_X2 U2135 ( .A(n271), .B(a[12]), .ZN(n2914) );
  AND3_X4 U2137 ( .A1(n2937), .A2(n2915), .A3(n2926), .ZN(n374) );
  XNOR2_X2 U2140 ( .A(n268), .B(a[9]), .ZN(n2915) );
  XNOR2_X2 U2145 ( .A(n265), .B(a[6]), .ZN(n2916) );
  AND3_X4 U2147 ( .A1(n2939), .A2(n2917), .A3(n2928), .ZN(n370) );
  XNOR2_X2 U2150 ( .A(n262), .B(a[3]), .ZN(n2917) );
  XOR2_X2 U2151 ( .A(a[4]), .B(n265), .Z(n2939) );
  AND3_X4 U2152 ( .A1(n2940), .A2(n2929), .A3(n2918), .ZN(n368) );
  XNOR2_X2 U2158 ( .A(n1441), .B(n1440), .ZN(n2843) );
  NAND2_X4 U2159 ( .A1(n1441), .A2(n484), .ZN(n2808) );
  XOR2_X2 U2162 ( .A(n1452), .B(n1407), .Z(n2844) );
  OAI21_X4 U2163 ( .B1(n1600), .B2(n1442), .A(n1443), .ZN(n1441) );
  NAND2_X4 U2164 ( .A1(n1528), .A2(n1444), .ZN(n1442) );
  AOI21_X4 U2165 ( .B1(n1529), .B2(n1444), .A(n1445), .ZN(n1443) );
  NOR2_X4 U2166 ( .A1(n1488), .A2(n1446), .ZN(n1444) );
  OAI21_X4 U2167 ( .B1(n1489), .B2(n1446), .A(n1447), .ZN(n1445) );
  NAND2_X4 U2168 ( .A1(n1468), .A2(n1448), .ZN(n1446) );
  AOI21_X4 U2169 ( .B1(n1448), .B2(n1469), .A(n1449), .ZN(n1447) );
  NOR2_X4 U2170 ( .A1(n1459), .A2(n1450), .ZN(n1448) );
  OAI21_X4 U2171 ( .B1(n1450), .B2(n1462), .A(n1451), .ZN(n1449) );
  NAND2_X4 U2172 ( .A1(n1689), .A2(n1451), .ZN(n1407) );
  NOR2_X4 U2174 ( .A1(n481), .A2(n484), .ZN(n1450) );
  NAND2_X4 U2175 ( .A1(n481), .A2(n484), .ZN(n1451) );
  XOR2_X2 U2176 ( .A(n1463), .B(n1408), .Z(n2845) );
  AOI21_X4 U2177 ( .B1(n1599), .B2(n1453), .A(n1454), .ZN(n1452) );
  NOR2_X4 U2178 ( .A1(n1530), .A2(n1455), .ZN(n1453) );
  OAI21_X4 U2179 ( .B1(n1531), .B2(n1455), .A(n1456), .ZN(n1454) );
  NAND2_X4 U2180 ( .A1(n1457), .A2(n1490), .ZN(n1455) );
  AOI21_X4 U2181 ( .B1(n1457), .B2(n1491), .A(n1458), .ZN(n1456) );
  NOR2_X4 U2182 ( .A1(n1470), .A2(n1459), .ZN(n1457) );
  OAI21_X4 U2183 ( .B1(n1471), .B2(n1459), .A(n1462), .ZN(n1458) );
  NAND2_X4 U2186 ( .A1(n1690), .A2(n1462), .ZN(n1408) );
  NOR2_X4 U2188 ( .A1(n478), .A2(n481), .ZN(n1459) );
  NAND2_X4 U2189 ( .A1(n478), .A2(n481), .ZN(n1462) );
  XOR2_X2 U2190 ( .A(n1476), .B(n1409), .Z(n2846) );
  AOI21_X4 U2191 ( .B1(n1599), .B2(n1464), .A(n1465), .ZN(n1463) );
  NOR2_X4 U2192 ( .A1(n1530), .A2(n1466), .ZN(n1464) );
  OAI21_X4 U2193 ( .B1(n1531), .B2(n1466), .A(n1467), .ZN(n1465) );
  NAND2_X4 U2194 ( .A1(n1490), .A2(n1468), .ZN(n1466) );
  AOI21_X4 U2195 ( .B1(n1491), .B2(n1468), .A(n1469), .ZN(n1467) );
  NOR2_X4 U2200 ( .A1(n1483), .A2(n1474), .ZN(n1468) );
  OAI21_X4 U2201 ( .B1(n1474), .B2(n1484), .A(n1475), .ZN(n1469) );
  NAND2_X4 U2202 ( .A1(n1691), .A2(n1475), .ZN(n1409) );
  NOR2_X4 U2204 ( .A1(n475), .A2(n478), .ZN(n1474) );
  NAND2_X4 U2205 ( .A1(n475), .A2(n478), .ZN(n1475) );
  XOR2_X2 U2206 ( .A(n1485), .B(n1410), .Z(n2847) );
  AOI21_X4 U2207 ( .B1(n1599), .B2(n1477), .A(n1478), .ZN(n1476) );
  NOR2_X4 U2208 ( .A1(n1530), .A2(n1479), .ZN(n1477) );
  OAI21_X4 U2209 ( .B1(n1531), .B2(n1479), .A(n1480), .ZN(n1478) );
  NAND2_X4 U2210 ( .A1(n1490), .A2(n1692), .ZN(n1479) );
  AOI21_X4 U2211 ( .B1(n1491), .B2(n1692), .A(n1482), .ZN(n1480) );
  NAND2_X4 U2214 ( .A1(n1692), .A2(n1484), .ZN(n1410) );
  NOR2_X4 U2216 ( .A1(n472), .A2(n475), .ZN(n1483) );
  NAND2_X4 U2217 ( .A1(n472), .A2(n475), .ZN(n1484) );
  XOR2_X2 U2218 ( .A(n1498), .B(n1411), .Z(n2848) );
  AOI21_X4 U2219 ( .B1(n1599), .B2(n1486), .A(n1487), .ZN(n1485) );
  NOR2_X4 U2220 ( .A1(n1530), .A2(n1488), .ZN(n1486) );
  OAI21_X4 U2221 ( .B1(n1531), .B2(n1488), .A(n1489), .ZN(n1487) );
  NAND2_X4 U2226 ( .A1(n1512), .A2(n1494), .ZN(n1488) );
  AOI21_X4 U2227 ( .B1(n1494), .B2(n1513), .A(n1495), .ZN(n1489) );
  NOR2_X4 U2228 ( .A1(n1505), .A2(n1496), .ZN(n1494) );
  OAI21_X4 U2229 ( .B1(n1496), .B2(n1506), .A(n1497), .ZN(n1495) );
  NAND2_X4 U2230 ( .A1(n1693), .A2(n1497), .ZN(n1411) );
  NOR2_X4 U2232 ( .A1(n469), .A2(n472), .ZN(n1496) );
  NAND2_X4 U2233 ( .A1(n469), .A2(n472), .ZN(n1497) );
  XOR2_X2 U2234 ( .A(n1507), .B(n1412), .Z(n2849) );
  AOI21_X4 U2235 ( .B1(n1599), .B2(n1499), .A(n1500), .ZN(n1498) );
  NOR2_X4 U2236 ( .A1(n1530), .A2(n1501), .ZN(n1499) );
  OAI21_X4 U2237 ( .B1(n1531), .B2(n1501), .A(n1502), .ZN(n1500) );
  NAND2_X4 U2238 ( .A1(n1512), .A2(n1694), .ZN(n1501) );
  AOI21_X4 U2239 ( .B1(n1513), .B2(n1694), .A(n1504), .ZN(n1502) );
  NAND2_X4 U2242 ( .A1(n1694), .A2(n1506), .ZN(n1412) );
  NOR2_X4 U2244 ( .A1(n466), .A2(n469), .ZN(n1505) );
  NAND2_X4 U2245 ( .A1(n466), .A2(n469), .ZN(n1506) );
  XOR2_X2 U2246 ( .A(n1520), .B(n1413), .Z(n2850) );
  AOI21_X4 U2247 ( .B1(n1599), .B2(n1508), .A(n1509), .ZN(n1507) );
  NOR2_X4 U2248 ( .A1(n1530), .A2(n1510), .ZN(n1508) );
  OAI21_X4 U2249 ( .B1(n1531), .B2(n1510), .A(n1511), .ZN(n1509) );
  NOR2_X4 U2256 ( .A1(n1523), .A2(n1518), .ZN(n1512) );
  OAI21_X4 U2257 ( .B1(n1518), .B2(n1526), .A(n1519), .ZN(n1513) );
  NAND2_X4 U2258 ( .A1(n1695), .A2(n1519), .ZN(n1413) );
  NOR2_X4 U2260 ( .A1(n463), .A2(n466), .ZN(n1518) );
  NAND2_X4 U2261 ( .A1(n463), .A2(n466), .ZN(n1519) );
  XOR2_X2 U2262 ( .A(n1527), .B(n1414), .Z(n2851) );
  AOI21_X4 U2263 ( .B1(n1599), .B2(n1521), .A(n1522), .ZN(n1520) );
  NOR2_X4 U2264 ( .A1(n1530), .A2(n1523), .ZN(n1521) );
  OAI21_X4 U2265 ( .B1(n1531), .B2(n1523), .A(n1526), .ZN(n1522) );
  NAND2_X4 U2268 ( .A1(n1696), .A2(n1526), .ZN(n1414) );
  NOR2_X4 U2270 ( .A1(n460), .A2(n463), .ZN(n1523) );
  NAND2_X4 U2271 ( .A1(n460), .A2(n463), .ZN(n1526) );
  XOR2_X2 U2272 ( .A(n1540), .B(n1415), .Z(n2852) );
  AOI21_X4 U2273 ( .B1(n1599), .B2(n1528), .A(n1529), .ZN(n1527) );
  NOR2_X4 U2278 ( .A1(n1568), .A2(n1534), .ZN(n1528) );
  OAI21_X4 U2279 ( .B1(n1569), .B2(n1534), .A(n1535), .ZN(n1529) );
  NAND2_X4 U2280 ( .A1(n1552), .A2(n1536), .ZN(n1534) );
  AOI21_X4 U2281 ( .B1(n1536), .B2(n1555), .A(n1537), .ZN(n1535) );
  NOR2_X4 U2282 ( .A1(n1543), .A2(n1538), .ZN(n1536) );
  OAI21_X4 U2283 ( .B1(n1538), .B2(n1546), .A(n1539), .ZN(n1537) );
  NAND2_X4 U2284 ( .A1(n1697), .A2(n1539), .ZN(n1415) );
  NOR2_X4 U2286 ( .A1(n457), .A2(n460), .ZN(n1538) );
  NAND2_X4 U2287 ( .A1(n457), .A2(n460), .ZN(n1539) );
  XOR2_X2 U2288 ( .A(n1547), .B(n1416), .Z(n2853) );
  AOI21_X4 U2289 ( .B1(n1599), .B2(n1541), .A(n1542), .ZN(n1540) );
  NOR2_X4 U2290 ( .A1(n1550), .A2(n1543), .ZN(n1541) );
  OAI21_X4 U2291 ( .B1(n1551), .B2(n1543), .A(n1546), .ZN(n1542) );
  NAND2_X4 U2294 ( .A1(n1698), .A2(n1546), .ZN(n1416) );
  NOR2_X4 U2296 ( .A1(n454), .A2(n457), .ZN(n1543) );
  NAND2_X4 U2297 ( .A1(n454), .A2(n457), .ZN(n1546) );
  XOR2_X2 U2298 ( .A(n1558), .B(n1417), .Z(n2854) );
  AOI21_X4 U2299 ( .B1(n1599), .B2(n1548), .A(n1549), .ZN(n1547) );
  NAND2_X4 U2302 ( .A1(n1570), .A2(n1552), .ZN(n1550) );
  AOI21_X4 U2303 ( .B1(n1571), .B2(n1552), .A(n1555), .ZN(n1551) );
  NOR2_X4 U2306 ( .A1(n1561), .A2(n1556), .ZN(n1552) );
  OAI21_X4 U2307 ( .B1(n1556), .B2(n1564), .A(n1557), .ZN(n1555) );
  NAND2_X4 U2308 ( .A1(n1699), .A2(n1557), .ZN(n1417) );
  NOR2_X4 U2310 ( .A1(n451), .A2(n454), .ZN(n1556) );
  NAND2_X4 U2311 ( .A1(n451), .A2(n454), .ZN(n1557) );
  XOR2_X2 U2312 ( .A(n1565), .B(n1418), .Z(n2855) );
  AOI21_X4 U2313 ( .B1(n1599), .B2(n1559), .A(n1560), .ZN(n1558) );
  NOR2_X4 U2314 ( .A1(n1568), .A2(n1561), .ZN(n1559) );
  OAI21_X4 U2315 ( .B1(n1569), .B2(n1561), .A(n1564), .ZN(n1560) );
  NAND2_X4 U2318 ( .A1(n1700), .A2(n1564), .ZN(n1418) );
  NOR2_X4 U2320 ( .A1(n448), .A2(n451), .ZN(n1561) );
  NAND2_X4 U2321 ( .A1(n448), .A2(n451), .ZN(n1564) );
  XOR2_X2 U2322 ( .A(n1578), .B(n1419), .Z(n2856) );
  AOI21_X4 U2323 ( .B1(n1599), .B2(n1570), .A(n1571), .ZN(n1565) );
  NAND2_X4 U2330 ( .A1(n1586), .A2(n1574), .ZN(n1568) );
  AOI21_X4 U2331 ( .B1(n1574), .B2(n1587), .A(n1575), .ZN(n1569) );
  NOR2_X4 U2332 ( .A1(n1581), .A2(n1576), .ZN(n1574) );
  OAI21_X4 U2333 ( .B1(n1576), .B2(n1584), .A(n1577), .ZN(n1575) );
  NAND2_X4 U2334 ( .A1(n1701), .A2(n1577), .ZN(n1419) );
  NOR2_X4 U2336 ( .A1(n445), .A2(n448), .ZN(n1576) );
  NAND2_X4 U2337 ( .A1(n445), .A2(n448), .ZN(n1577) );
  XOR2_X2 U2338 ( .A(n1585), .B(n1420), .Z(n2857) );
  AOI21_X4 U2339 ( .B1(n1599), .B2(n1579), .A(n1580), .ZN(n1578) );
  NOR2_X4 U2340 ( .A1(n1588), .A2(n1581), .ZN(n1579) );
  OAI21_X4 U2341 ( .B1(n1589), .B2(n1581), .A(n1584), .ZN(n1580) );
  NAND2_X4 U2344 ( .A1(n1702), .A2(n1584), .ZN(n1420) );
  NOR2_X4 U2346 ( .A1(n442), .A2(n445), .ZN(n1581) );
  NAND2_X4 U2347 ( .A1(n442), .A2(n445), .ZN(n1584) );
  XOR2_X2 U2348 ( .A(n1594), .B(n1421), .Z(n2858) );
  AOI21_X4 U2349 ( .B1(n1599), .B2(n1586), .A(n1587), .ZN(n1585) );
  NOR2_X4 U2354 ( .A1(n1597), .A2(n1592), .ZN(n1586) );
  OAI21_X4 U2355 ( .B1(n1592), .B2(n1598), .A(n1593), .ZN(n1587) );
  NAND2_X4 U2356 ( .A1(n1703), .A2(n1593), .ZN(n1421) );
  NOR2_X4 U2358 ( .A1(n439), .A2(n442), .ZN(n1592) );
  NAND2_X4 U2359 ( .A1(n439), .A2(n442), .ZN(n1593) );
  XNOR2_X2 U2360 ( .A(n1599), .B(n1422), .ZN(n2859) );
  AOI21_X4 U2361 ( .B1(n1599), .B2(n1704), .A(n1596), .ZN(n1594) );
  NAND2_X4 U2364 ( .A1(n1704), .A2(n1598), .ZN(n1422) );
  NOR2_X4 U2366 ( .A1(n436), .A2(n439), .ZN(n1597) );
  NAND2_X4 U2367 ( .A1(n436), .A2(n439), .ZN(n1598) );
  XOR2_X2 U2368 ( .A(n1609), .B(n1423), .Z(n2860) );
  AOI21_X4 U2370 ( .B1(n1655), .B2(n1601), .A(n1602), .ZN(n1600) );
  NOR2_X4 U2371 ( .A1(n1629), .A2(n1603), .ZN(n1601) );
  OAI21_X4 U2372 ( .B1(n1630), .B2(n1603), .A(n1604), .ZN(n1602) );
  NAND2_X4 U2373 ( .A1(n1617), .A2(n1605), .ZN(n1603) );
  AOI21_X4 U2374 ( .B1(n1605), .B2(n1620), .A(n1606), .ZN(n1604) );
  NOR2_X4 U2375 ( .A1(n1612), .A2(n1607), .ZN(n1605) );
  OAI21_X4 U2376 ( .B1(n1607), .B2(n1613), .A(n1608), .ZN(n1606) );
  NAND2_X4 U2377 ( .A1(n1705), .A2(n1608), .ZN(n1423) );
  NOR2_X4 U2379 ( .A1(n433), .A2(n436), .ZN(n1607) );
  NAND2_X4 U2380 ( .A1(n433), .A2(n436), .ZN(n1608) );
  XNOR2_X2 U2381 ( .A(n1614), .B(n1424), .ZN(n2861) );
  AOI21_X4 U2382 ( .B1(n1614), .B2(n1706), .A(n1611), .ZN(n1609) );
  NAND2_X4 U2385 ( .A1(n1706), .A2(n1613), .ZN(n1424) );
  NOR2_X4 U2387 ( .A1(n430), .A2(n433), .ZN(n1612) );
  NAND2_X4 U2388 ( .A1(n430), .A2(n433), .ZN(n1613) );
  XOR2_X2 U2389 ( .A(n1623), .B(n1425), .Z(n2862) );
  OAI21_X4 U2390 ( .B1(n1654), .B2(n1615), .A(n1616), .ZN(n1614) );
  NAND2_X4 U2391 ( .A1(n1631), .A2(n1617), .ZN(n1615) );
  AOI21_X4 U2392 ( .B1(n1632), .B2(n1617), .A(n1620), .ZN(n1616) );
  NOR2_X4 U2395 ( .A1(n1626), .A2(n1621), .ZN(n1617) );
  OAI21_X4 U2396 ( .B1(n1621), .B2(n1627), .A(n1622), .ZN(n1620) );
  NAND2_X4 U2397 ( .A1(n1707), .A2(n1622), .ZN(n1425) );
  NOR2_X4 U2399 ( .A1(n427), .A2(n430), .ZN(n1621) );
  NAND2_X4 U2400 ( .A1(n427), .A2(n430), .ZN(n1622) );
  XNOR2_X2 U2401 ( .A(n1628), .B(n1426), .ZN(n2863) );
  AOI21_X4 U2402 ( .B1(n1628), .B2(n1708), .A(n1625), .ZN(n1623) );
  NAND2_X4 U2405 ( .A1(n1708), .A2(n1627), .ZN(n1426) );
  NOR2_X4 U2407 ( .A1(n424), .A2(n427), .ZN(n1626) );
  NAND2_X4 U2408 ( .A1(n424), .A2(n427), .ZN(n1627) );
  XOR2_X2 U2409 ( .A(n1639), .B(n1427), .Z(n2864) );
  OAI21_X4 U2410 ( .B1(n1654), .B2(n1629), .A(n1630), .ZN(n1628) );
  NAND2_X4 U2415 ( .A1(n1647), .A2(n1635), .ZN(n1629) );
  AOI21_X4 U2416 ( .B1(n1635), .B2(n1648), .A(n1636), .ZN(n1630) );
  NOR2_X4 U2417 ( .A1(n1642), .A2(n1637), .ZN(n1635) );
  OAI21_X4 U2418 ( .B1(n1637), .B2(n1643), .A(n1638), .ZN(n1636) );
  NAND2_X4 U2419 ( .A1(n1709), .A2(n1638), .ZN(n1427) );
  NOR2_X4 U2421 ( .A1(n421), .A2(n424), .ZN(n1637) );
  NAND2_X4 U2422 ( .A1(n421), .A2(n424), .ZN(n1638) );
  XNOR2_X2 U2423 ( .A(n1644), .B(n1428), .ZN(n2865) );
  AOI21_X4 U2424 ( .B1(n1644), .B2(n1710), .A(n1641), .ZN(n1639) );
  NAND2_X4 U2427 ( .A1(n1710), .A2(n1643), .ZN(n1428) );
  NOR2_X4 U2429 ( .A1(n418), .A2(n421), .ZN(n1642) );
  NAND2_X4 U2430 ( .A1(n418), .A2(n421), .ZN(n1643) );
  XNOR2_X2 U2431 ( .A(n1651), .B(n1429), .ZN(n2866) );
  OAI21_X4 U2432 ( .B1(n1654), .B2(n1645), .A(n1646), .ZN(n1644) );
  NOR2_X4 U2435 ( .A1(n1652), .A2(n1649), .ZN(n1647) );
  OAI21_X4 U2436 ( .B1(n1649), .B2(n1653), .A(n1650), .ZN(n1648) );
  NAND2_X4 U2437 ( .A1(n1711), .A2(n1650), .ZN(n1429) );
  NOR2_X4 U2439 ( .A1(n415), .A2(n418), .ZN(n1649) );
  NAND2_X4 U2440 ( .A1(n415), .A2(n418), .ZN(n1650) );
  XOR2_X2 U2441 ( .A(n1654), .B(n1430), .Z(n2867) );
  OAI21_X4 U2442 ( .B1(n1654), .B2(n1652), .A(n1653), .ZN(n1651) );
  NAND2_X4 U2443 ( .A1(n1712), .A2(n1653), .ZN(n1430) );
  NOR2_X4 U2445 ( .A1(n412), .A2(n415), .ZN(n1652) );
  NAND2_X4 U2446 ( .A1(n412), .A2(n415), .ZN(n1653) );
  XNOR2_X2 U2447 ( .A(n1662), .B(n1431), .ZN(n2868) );
  OAI21_X4 U2449 ( .B1(n1676), .B2(n1656), .A(n1657), .ZN(n1655) );
  NAND2_X4 U2450 ( .A1(n1666), .A2(n1658), .ZN(n1656) );
  AOI21_X4 U2451 ( .B1(n1658), .B2(n1667), .A(n1659), .ZN(n1657) );
  NOR2_X4 U2452 ( .A1(n1663), .A2(n1660), .ZN(n1658) );
  OAI21_X4 U2453 ( .B1(n1660), .B2(n1664), .A(n1661), .ZN(n1659) );
  NAND2_X4 U2454 ( .A1(n1713), .A2(n1661), .ZN(n1431) );
  NOR2_X4 U2456 ( .A1(n409), .A2(n412), .ZN(n1660) );
  NAND2_X4 U2457 ( .A1(n409), .A2(n412), .ZN(n1661) );
  XOR2_X2 U2458 ( .A(n1665), .B(n1432), .Z(n2869) );
  OAI21_X4 U2459 ( .B1(n1665), .B2(n1663), .A(n1664), .ZN(n1662) );
  NAND2_X4 U2460 ( .A1(n1714), .A2(n1664), .ZN(n1432) );
  NOR2_X4 U2462 ( .A1(n406), .A2(n409), .ZN(n1663) );
  NAND2_X4 U2463 ( .A1(n406), .A2(n409), .ZN(n1664) );
  XOR2_X2 U2464 ( .A(n1670), .B(n1433), .Z(n2870) );
  AOI21_X4 U2465 ( .B1(n1675), .B2(n1666), .A(n1667), .ZN(n1665) );
  NOR2_X4 U2466 ( .A1(n1673), .A2(n1668), .ZN(n1666) );
  OAI21_X4 U2467 ( .B1(n1668), .B2(n1674), .A(n1669), .ZN(n1667) );
  NAND2_X4 U2468 ( .A1(n1715), .A2(n1669), .ZN(n1433) );
  NOR2_X4 U2470 ( .A1(n403), .A2(n406), .ZN(n1668) );
  NAND2_X4 U2471 ( .A1(n403), .A2(n406), .ZN(n1669) );
  XNOR2_X2 U2472 ( .A(n1675), .B(n1434), .ZN(n2871) );
  AOI21_X4 U2473 ( .B1(n1675), .B2(n1716), .A(n1672), .ZN(n1670) );
  NAND2_X4 U2476 ( .A1(n1716), .A2(n1674), .ZN(n1434) );
  NOR2_X4 U2478 ( .A1(n400), .A2(n403), .ZN(n1673) );
  NAND2_X4 U2479 ( .A1(n400), .A2(n403), .ZN(n1674) );
  XNOR2_X2 U2480 ( .A(n1681), .B(n1435), .ZN(n2872) );
  AOI21_X4 U2482 ( .B1(n1677), .B2(n1685), .A(n1678), .ZN(n1676) );
  NOR2_X4 U2483 ( .A1(n1682), .A2(n1679), .ZN(n1677) );
  OAI21_X4 U2484 ( .B1(n1679), .B2(n1683), .A(n1680), .ZN(n1678) );
  NAND2_X4 U2485 ( .A1(n1717), .A2(n1680), .ZN(n1435) );
  NOR2_X4 U2487 ( .A1(n397), .A2(n400), .ZN(n1679) );
  NAND2_X4 U2488 ( .A1(n397), .A2(n400), .ZN(n1680) );
  XOR2_X2 U2489 ( .A(n1436), .B(n1684), .Z(n2873) );
  OAI21_X4 U2490 ( .B1(n1682), .B2(n1684), .A(n1683), .ZN(n1681) );
  NAND2_X4 U2491 ( .A1(n1718), .A2(n1683), .ZN(n1436) );
  NOR2_X4 U2493 ( .A1(n393), .A2(n397), .ZN(n1682) );
  NAND2_X4 U2494 ( .A1(n393), .A2(n397), .ZN(n1683) );
  NAND2_X4 U2498 ( .A1(n1719), .A2(n1684), .ZN(n2840) );
  NOR2_X4 U2500 ( .A1(n390), .A2(n393), .ZN(n1686) );
  NAND2_X4 U2501 ( .A1(n390), .A2(n393), .ZN(n1684) );
  INV_X1 U2506 ( .A(n271), .ZN(n3220) );
  XNOR2_X1 U2507 ( .A(n280), .B(a[21]), .ZN(n2911) );
  XOR2_X1 U2508 ( .A(a[22]), .B(n283), .Z(n2933) );
  XNOR2_X1 U2509 ( .A(a[21]), .B(a[22]), .ZN(n2922) );
  XNOR2_X1 U2510 ( .A(n283), .B(a[24]), .ZN(n2910) );
  XOR2_X1 U2511 ( .A(a[25]), .B(n286), .Z(n2932) );
  XNOR2_X1 U2512 ( .A(a[24]), .B(a[25]), .ZN(n2921) );
  XOR2_X1 U2513 ( .A(a[28]), .B(n289), .Z(n2931) );
  XNOR2_X1 U2514 ( .A(a[27]), .B(a[28]), .ZN(n2920) );
  XOR2_X1 U2515 ( .A(a[1]), .B(n262), .Z(n2940) );
  XNOR2_X1 U2516 ( .A(a[3]), .B(a[4]), .ZN(n2928) );
  XNOR2_X1 U2517 ( .A(a[6]), .B(a[7]), .ZN(n2927) );
  INV_X1 U2518 ( .A(a[10]), .ZN(n3222) );
  XNOR2_X1 U2519 ( .A(a[9]), .B(a[10]), .ZN(n2926) );
  XOR2_X1 U2520 ( .A(a[13]), .B(n274), .Z(n2936) );
  XNOR2_X1 U2521 ( .A(a[12]), .B(a[13]), .ZN(n2925) );
  XNOR2_X1 U2522 ( .A(n274), .B(a[15]), .ZN(n2913) );
  XOR2_X1 U2523 ( .A(a[16]), .B(n277), .Z(n2935) );
  XNOR2_X1 U2524 ( .A(a[15]), .B(a[16]), .ZN(n2924) );
  XNOR2_X1 U2525 ( .A(n277), .B(a[18]), .ZN(n2912) );
  XOR2_X1 U2526 ( .A(a[19]), .B(n280), .Z(n2934) );
  XNOR2_X1 U2527 ( .A(a[18]), .B(a[19]), .ZN(n2923) );
  XNOR2_X1 U2528 ( .A(a[0]), .B(a[1]), .ZN(n2929) );
  OR2_X1 U2529 ( .A1(n2929), .A2(a[0]), .ZN(n3238) );
  INV_X1 U2530 ( .A(a[0]), .ZN(n2918) );
  XNOR2_X1 U2531 ( .A(a[30]), .B(a[31]), .ZN(n2919) );
  NAND3_X1 U2532 ( .A1(n2938), .A2(n2916), .A3(n2927), .ZN(n3126) );
  INV_X1 U2533 ( .A(n3126), .ZN(n3127) );
  INV_X1 U2534 ( .A(n3126), .ZN(n3128) );
  BUF_X1 U2535 ( .A(n354), .Z(n3129) );
  BUF_X1 U2536 ( .A(n351), .Z(n3130) );
  BUF_X1 U2537 ( .A(n348), .Z(n3131) );
  INV_X1 U2538 ( .A(n2914), .ZN(n3234) );
  BUF_X1 U2539 ( .A(n345), .Z(n3132) );
  BUF_X1 U2540 ( .A(n336), .Z(n3133) );
  OR2_X1 U2541 ( .A1(n2933), .A2(n2911), .ZN(n3134) );
  INV_X1 U2542 ( .A(n3134), .ZN(n3135) );
  INV_X1 U2543 ( .A(n3134), .ZN(n3136) );
  OR2_X1 U2544 ( .A1(n2934), .A2(n2912), .ZN(n3137) );
  INV_X1 U2545 ( .A(n3137), .ZN(n3138) );
  INV_X1 U2546 ( .A(n3137), .ZN(n3139) );
  OR2_X1 U2547 ( .A1(n2935), .A2(n2913), .ZN(n3140) );
  INV_X1 U2548 ( .A(n3140), .ZN(n3141) );
  INV_X1 U2549 ( .A(n3140), .ZN(n3142) );
  OR2_X1 U2550 ( .A1(n2908), .A2(a[31]), .ZN(n3143) );
  INV_X1 U2551 ( .A(n3143), .ZN(n3144) );
  INV_X1 U2552 ( .A(n3143), .ZN(n3145) );
  XNOR2_X1 U2553 ( .A(n289), .B(a[30]), .ZN(n2908) );
  OR2_X1 U2554 ( .A1(n2931), .A2(n2909), .ZN(n3146) );
  INV_X1 U2555 ( .A(n3146), .ZN(n3147) );
  INV_X1 U2556 ( .A(n3146), .ZN(n3148) );
  XNOR2_X1 U2557 ( .A(n286), .B(a[27]), .ZN(n2909) );
  OR2_X1 U2558 ( .A1(n2932), .A2(n2910), .ZN(n3149) );
  INV_X1 U2559 ( .A(n3149), .ZN(n3150) );
  INV_X1 U2560 ( .A(n3149), .ZN(n3151) );
  OR2_X1 U2561 ( .A1(n2940), .A2(n2918), .ZN(n3152) );
  INV_X1 U2562 ( .A(n3152), .ZN(n3153) );
  INV_X1 U2563 ( .A(n3152), .ZN(n3154) );
  AND2_X1 U2564 ( .A1(a[31]), .A2(n3228), .ZN(n3155) );
  INV_X1 U2565 ( .A(n3155), .ZN(n3156) );
  INV_X4 U2566 ( .A(n3155), .ZN(n3157) );
  AND2_X1 U2567 ( .A1(n2931), .A2(n3229), .ZN(n3158) );
  INV_X1 U2568 ( .A(n3158), .ZN(n3159) );
  INV_X4 U2569 ( .A(n3158), .ZN(n3160) );
  BUF_X1 U2570 ( .A(n360), .Z(n3161) );
  NAND2_X4 U2571 ( .A1(n2932), .A2(n3230), .ZN(n360) );
  BUF_X1 U2572 ( .A(n357), .Z(n3162) );
  NAND2_X4 U2573 ( .A1(n2933), .A2(n3231), .ZN(n357) );
  XOR2_X1 U2574 ( .A(n719), .B(n718), .Z(n3163) );
  XOR2_X1 U2575 ( .A(n520), .B(n3163), .Z(product[62]) );
  NAND2_X1 U2576 ( .A1(n520), .A2(n719), .ZN(n3164) );
  NAND2_X1 U2577 ( .A1(n520), .A2(n718), .ZN(n3165) );
  NAND2_X1 U2578 ( .A1(n719), .A2(n718), .ZN(n3166) );
  NAND3_X1 U2579 ( .A1(n3164), .A2(n3166), .A3(n3165), .ZN(n519) );
  BUF_X1 U2580 ( .A(n524), .Z(n3167) );
  BUF_X1 U2581 ( .A(n534), .Z(n3168) );
  XOR2_X1 U2582 ( .A(n743), .B(n739), .Z(n3169) );
  XOR2_X1 U2583 ( .A(n526), .B(n3169), .Z(product[56]) );
  NAND2_X1 U2584 ( .A1(n526), .A2(n743), .ZN(n3170) );
  NAND2_X1 U2585 ( .A1(n526), .A2(n739), .ZN(n3171) );
  NAND2_X1 U2586 ( .A1(n743), .A2(n739), .ZN(n3172) );
  NAND3_X2 U2587 ( .A1(n3170), .A2(n3172), .A3(n3171), .ZN(n525) );
  XOR2_X1 U2588 ( .A(n825), .B(n836), .Z(n3173) );
  XOR2_X1 U2589 ( .A(n536), .B(n3173), .Z(product[46]) );
  NAND2_X1 U2590 ( .A1(n536), .A2(n825), .ZN(n3174) );
  NAND2_X1 U2591 ( .A1(n536), .A2(n836), .ZN(n3175) );
  NAND2_X1 U2592 ( .A1(n825), .A2(n836), .ZN(n3176) );
  NAND3_X2 U2593 ( .A1(n3174), .A2(n3176), .A3(n3175), .ZN(n535) );
  XOR2_X1 U2594 ( .A(n996), .B(n979), .Z(n3177) );
  XOR2_X1 U2595 ( .A(n546), .B(n3177), .Z(product[36]) );
  NAND2_X1 U2596 ( .A1(n546), .A2(n996), .ZN(n3178) );
  NAND2_X1 U2597 ( .A1(n546), .A2(n979), .ZN(n3179) );
  NAND2_X1 U2598 ( .A1(n996), .A2(n979), .ZN(n3180) );
  NAND3_X2 U2599 ( .A1(n3178), .A2(n3180), .A3(n3179), .ZN(n545) );
  BUF_X1 U2600 ( .A(n555), .Z(n3181) );
  BUF_X1 U2601 ( .A(n619), .Z(n3182) );
  BUF_X1 U2602 ( .A(n635), .Z(n3183) );
  INV_X1 U2603 ( .A(n717), .ZN(n718) );
  NAND3_X1 U2604 ( .A1(n3187), .A2(n3188), .A3(n3189), .ZN(n524) );
  NAND3_X1 U2605 ( .A1(n3195), .A2(n3196), .A3(n3197), .ZN(n534) );
  OAI21_X1 U2606 ( .B1(n558), .B2(n556), .A(n557), .ZN(n555) );
  AOI21_X4 U2607 ( .B1(n571), .B2(n688), .A(n568), .ZN(n566) );
  OAI21_X1 U2608 ( .B1(n638), .B2(n636), .A(n637), .ZN(n635) );
  XNOR2_X1 U2609 ( .A(n515), .B(n667), .ZN(product[5]) );
  XOR2_X2 U2610 ( .A(a[7]), .B(n268), .Z(n2938) );
  OAI21_X1 U2611 ( .B1(n2839), .B2(n342), .A(n2669), .ZN(n2635) );
  AOI222_X1 U2612 ( .A1(n295), .A2(n397), .B1(n317), .B2(n393), .C1(n3127), 
        .C2(n390), .ZN(n2669) );
  INV_X1 U2613 ( .A(n299), .ZN(n3184) );
  INV_X4 U2614 ( .A(n3184), .ZN(n3185) );
  NOR2_X2 U2615 ( .A1(n2936), .A2(n2914), .ZN(n299) );
  OAI21_X2 U2616 ( .B1(n670), .B2(n668), .A(n669), .ZN(n667) );
  XNOR2_X1 U2617 ( .A(n3183), .B(n507), .ZN(product[13]) );
  XOR2_X1 U2618 ( .A(n638), .B(n508), .Z(product[12]) );
  AOI21_X2 U2619 ( .B1(n643), .B2(n706), .A(n640), .ZN(n638) );
  XNOR2_X1 U2620 ( .A(n627), .B(n505), .ZN(product[15]) );
  XOR2_X1 U2621 ( .A(n630), .B(n506), .Z(product[14]) );
  OAI21_X2 U2622 ( .B1(n630), .B2(n628), .A(n629), .ZN(n627) );
  XOR2_X1 U2623 ( .A(n738), .B(n733), .Z(n3186) );
  XOR2_X1 U2624 ( .A(n3186), .B(n525), .Z(product[57]) );
  NAND2_X2 U2625 ( .A1(n738), .A2(n733), .ZN(n3187) );
  NAND2_X1 U2626 ( .A1(n738), .A2(n525), .ZN(n3188) );
  NAND2_X1 U2627 ( .A1(n733), .A2(n525), .ZN(n3189) );
  XOR2_X1 U2628 ( .A(n729), .B(n732), .Z(n3190) );
  XOR2_X1 U2629 ( .A(n3190), .B(n3167), .Z(product[58]) );
  NAND2_X1 U2630 ( .A1(n729), .A2(n732), .ZN(n3191) );
  NAND2_X1 U2631 ( .A1(n729), .A2(n524), .ZN(n3192) );
  NAND2_X1 U2632 ( .A1(n732), .A2(n524), .ZN(n3193) );
  NAND3_X1 U2633 ( .A1(n3191), .A2(n3192), .A3(n3193), .ZN(n523) );
  XOR2_X1 U2634 ( .A(n814), .B(n824), .Z(n3194) );
  XOR2_X1 U2635 ( .A(n3194), .B(n535), .Z(product[47]) );
  NAND2_X2 U2636 ( .A1(n814), .A2(n824), .ZN(n3195) );
  NAND2_X1 U2637 ( .A1(n814), .A2(n535), .ZN(n3196) );
  NAND2_X1 U2638 ( .A1(n824), .A2(n535), .ZN(n3197) );
  XOR2_X1 U2639 ( .A(n802), .B(n813), .Z(n3198) );
  XOR2_X1 U2640 ( .A(n3198), .B(n3168), .Z(product[48]) );
  NAND2_X1 U2641 ( .A1(n802), .A2(n813), .ZN(n3199) );
  NAND2_X1 U2642 ( .A1(n802), .A2(n534), .ZN(n3200) );
  NAND2_X1 U2643 ( .A1(n813), .A2(n534), .ZN(n3201) );
  NAND3_X1 U2644 ( .A1(n3199), .A2(n3200), .A3(n3201), .ZN(n533) );
  XOR2_X1 U2645 ( .A(n961), .B(n978), .Z(n3202) );
  XOR2_X1 U2646 ( .A(n3202), .B(n545), .Z(product[37]) );
  NAND2_X2 U2647 ( .A1(n961), .A2(n978), .ZN(n3203) );
  NAND2_X1 U2648 ( .A1(n961), .A2(n545), .ZN(n3204) );
  NAND2_X1 U2649 ( .A1(n978), .A2(n545), .ZN(n3205) );
  NAND3_X2 U2650 ( .A1(n3203), .A2(n3204), .A3(n3205), .ZN(n544) );
  XOR2_X1 U2651 ( .A(n944), .B(n960), .Z(n3206) );
  XOR2_X1 U2652 ( .A(n3206), .B(n544), .Z(product[38]) );
  NAND2_X1 U2653 ( .A1(n944), .A2(n960), .ZN(n3207) );
  NAND2_X1 U2654 ( .A1(n944), .A2(n544), .ZN(n3208) );
  NAND2_X1 U2655 ( .A1(n960), .A2(n544), .ZN(n3209) );
  NAND3_X1 U2656 ( .A1(n3207), .A2(n3208), .A3(n3209), .ZN(n543) );
  NAND2_X1 U2657 ( .A1(n519), .A2(n3223), .ZN(n3212) );
  NAND2_X1 U2658 ( .A1(n3210), .A2(n3211), .ZN(n3213) );
  NAND2_X1 U2659 ( .A1(n3212), .A2(n3213), .ZN(product[63]) );
  INV_X1 U2660 ( .A(n519), .ZN(n3210) );
  INV_X1 U2661 ( .A(n3223), .ZN(n3211) );
  BUF_X1 U2662 ( .A(n571), .Z(n3214) );
  BUF_X1 U2663 ( .A(n563), .Z(n3215) );
  BUF_X1 U2664 ( .A(n611), .Z(n3216) );
  BUF_X1 U2665 ( .A(n579), .Z(n3217) );
  BUF_X1 U2666 ( .A(n651), .Z(n3218) );
  BUF_X1 U2667 ( .A(n643), .Z(n3219) );
  INV_X1 U2668 ( .A(n485), .ZN(n3223) );
  OAI21_X1 U2669 ( .B1(n644), .B2(n646), .A(n645), .ZN(n643) );
  OAI21_X1 U2670 ( .B1(n2840), .B2(n342), .A(n2670), .ZN(n2636) );
  NAND2_X1 U2671 ( .A1(n715), .A2(n682), .ZN(n518) );
  NOR2_X1 U2672 ( .A1(n2093), .A2(n262), .ZN(n681) );
  NAND2_X2 U2673 ( .A1(n2093), .A2(n262), .ZN(n682) );
  NAND2_X4 U2674 ( .A1(n2934), .A2(n3232), .ZN(n354) );
  OR2_X4 U2675 ( .A1(n2926), .A2(n3235), .ZN(n3241) );
  INV_X8 U2676 ( .A(n3241), .ZN(n319) );
  XNOR2_X2 U2677 ( .A(n2569), .B(n3220), .ZN(n1988) );
  OR2_X4 U2678 ( .A1(n2939), .A2(n2917), .ZN(n3221) );
  INV_X32 U2679 ( .A(n3221), .ZN(n293) );
  NOR2_X1 U2680 ( .A1(n1351), .A2(n1356), .ZN(n649) );
  NAND2_X2 U2681 ( .A1(n1351), .A2(n1356), .ZN(n650) );
  XNOR2_X2 U2682 ( .A(n3222), .B(n271), .ZN(n2937) );
  NOR2_X2 U2683 ( .A1(n2090), .A2(n1373), .ZN(n673) );
  NAND2_X2 U2684 ( .A1(n1373), .A2(n2090), .ZN(n674) );
  AOI22_X1 U2685 ( .A1(n293), .A2(n393), .B1(n315), .B2(n390), .ZN(n2738) );
  OAI21_X1 U2686 ( .B1(n2840), .B2(n339), .A(n2738), .ZN(n2704) );
  INV_X8 U2687 ( .A(n3239), .ZN(n315) );
  OR2_X4 U2688 ( .A1(n2937), .A2(n2915), .ZN(n3224) );
  INV_X32 U2689 ( .A(n3224), .ZN(n297) );
  INV_X8 U2690 ( .A(n3240), .ZN(n317) );
  XNOR2_X2 U2691 ( .A(n2705), .B(n3225), .ZN(n2058) );
  INV_X32 U2692 ( .A(n265), .ZN(n3225) );
  NAND2_X4 U2693 ( .A1(n2935), .A2(n3233), .ZN(n351) );
  XNOR2_X1 U2694 ( .A(n3218), .B(n511), .ZN(product[9]) );
  XNOR2_X1 U2695 ( .A(n513), .B(n659), .ZN(product[7]) );
  OR2_X4 U2696 ( .A1(n2938), .A2(n2916), .ZN(n3226) );
  INV_X32 U2697 ( .A(n3226), .ZN(n295) );
  XNOR2_X1 U2698 ( .A(n2637), .B(n3227), .ZN(n2023) );
  INV_X32 U2699 ( .A(n268), .ZN(n3227) );
  AOI21_X4 U2700 ( .B1(n651), .B2(n708), .A(n648), .ZN(n646) );
  XOR2_X1 U2701 ( .A(n550), .B(n486), .Z(product[34]) );
  OAI21_X1 U2702 ( .B1(n550), .B2(n548), .A(n549), .ZN(n547) );
  AOI21_X2 U2703 ( .B1(n555), .B2(n684), .A(n552), .ZN(n550) );
  NAND2_X4 U2704 ( .A1(n2936), .A2(n3234), .ZN(n348) );
  NAND2_X4 U2705 ( .A1(n2940), .A2(a[0]), .ZN(n336) );
  NAND2_X4 U2706 ( .A1(n2937), .A2(n3235), .ZN(n345) );
  XNOR2_X1 U2707 ( .A(n3215), .B(n489), .ZN(product[31]) );
  XNOR2_X1 U2708 ( .A(n3181), .B(n487), .ZN(product[33]) );
  XNOR2_X1 U2709 ( .A(n3219), .B(n509), .ZN(product[11]) );
  NAND2_X4 U2710 ( .A1(n2938), .A2(n3236), .ZN(n342) );
  OAI21_X1 U2711 ( .B1(n2841), .B2(n342), .A(n2671), .ZN(n2637) );
  XNOR2_X1 U2712 ( .A(n3217), .B(n493), .ZN(product[27]) );
  XNOR2_X1 U2713 ( .A(n3182), .B(n503), .ZN(product[17]) );
  XNOR2_X1 U2714 ( .A(n3214), .B(n491), .ZN(product[29]) );
  XNOR2_X1 U2715 ( .A(n3216), .B(n501), .ZN(product[19]) );
  XOR2_X1 U2716 ( .A(n566), .B(n490), .Z(product[30]) );
  XOR2_X1 U2717 ( .A(n510), .B(n646), .Z(product[10]) );
  OAI21_X2 U2718 ( .B1(n566), .B2(n564), .A(n565), .ZN(n563) );
  NAND2_X4 U2719 ( .A1(n2939), .A2(n3237), .ZN(n339) );
  OAI21_X2 U2720 ( .B1(n654), .B2(n652), .A(n653), .ZN(n651) );
  OAI21_X2 U2721 ( .B1(n660), .B2(n662), .A(n661), .ZN(n659) );
  OAI21_X2 U2722 ( .B1(n614), .B2(n612), .A(n613), .ZN(n611) );
  OAI21_X2 U2723 ( .B1(n582), .B2(n580), .A(n581), .ZN(n579) );
  OAI21_X2 U2724 ( .B1(n574), .B2(n572), .A(n573), .ZN(n571) );
  OAI21_X2 U2725 ( .B1(n622), .B2(n620), .A(n621), .ZN(n619) );
  INV_X2 U2726 ( .A(n518), .ZN(product[0]) );
  INV_X2 U2727 ( .A(n941), .ZN(n959) );
  INV_X2 U2728 ( .A(n907), .ZN(n908) );
  INV_X2 U2729 ( .A(n891), .ZN(n892) );
  INV_X2 U2730 ( .A(n848), .ZN(n862) );
  INV_X2 U2731 ( .A(n811), .ZN(n823) );
  INV_X2 U2732 ( .A(n780), .ZN(n790) );
  INV_X2 U2733 ( .A(n755), .ZN(n763) );
  INV_X2 U2734 ( .A(n736), .ZN(n742) );
  INV_X2 U2735 ( .A(n723), .ZN(n727) );
  INV_X2 U2736 ( .A(n1720), .ZN(n716) );
  INV_X2 U2737 ( .A(n681), .ZN(n715) );
  INV_X2 U2738 ( .A(n668), .ZN(n713) );
  INV_X2 U2739 ( .A(n660), .ZN(n711) );
  INV_X2 U2740 ( .A(n652), .ZN(n709) );
  INV_X2 U2741 ( .A(n644), .ZN(n707) );
  INV_X2 U2742 ( .A(n636), .ZN(n705) );
  INV_X2 U2743 ( .A(n628), .ZN(n703) );
  INV_X2 U2744 ( .A(n620), .ZN(n701) );
  INV_X2 U2745 ( .A(n612), .ZN(n699) );
  INV_X2 U2746 ( .A(n604), .ZN(n697) );
  INV_X2 U2747 ( .A(n596), .ZN(n695) );
  INV_X2 U2748 ( .A(n588), .ZN(n693) );
  INV_X2 U2749 ( .A(n580), .ZN(n691) );
  INV_X2 U2750 ( .A(n572), .ZN(n689) );
  INV_X2 U2751 ( .A(n564), .ZN(n687) );
  INV_X2 U2752 ( .A(n556), .ZN(n685) );
  INV_X2 U2753 ( .A(n548), .ZN(n683) );
  INV_X2 U2754 ( .A(n682), .ZN(n680) );
  INV_X2 U2755 ( .A(n678), .ZN(n679) );
  INV_X2 U2756 ( .A(n2091), .ZN(n676) );
  INV_X2 U2757 ( .A(n674), .ZN(n672) );
  INV_X2 U2758 ( .A(n673), .ZN(n714) );
  INV_X2 U2759 ( .A(n666), .ZN(n664) );
  INV_X2 U2760 ( .A(n665), .ZN(n712) );
  INV_X2 U2761 ( .A(n658), .ZN(n656) );
  INV_X2 U2762 ( .A(n657), .ZN(n710) );
  INV_X2 U2763 ( .A(n650), .ZN(n648) );
  INV_X2 U2764 ( .A(n649), .ZN(n708) );
  INV_X2 U2765 ( .A(n642), .ZN(n640) );
  INV_X2 U2766 ( .A(n641), .ZN(n706) );
  INV_X2 U2767 ( .A(n634), .ZN(n632) );
  INV_X2 U2768 ( .A(n633), .ZN(n704) );
  INV_X2 U2769 ( .A(n626), .ZN(n624) );
  INV_X2 U2770 ( .A(n625), .ZN(n702) );
  INV_X2 U2771 ( .A(n618), .ZN(n616) );
  INV_X2 U2772 ( .A(n617), .ZN(n700) );
  INV_X2 U2773 ( .A(n610), .ZN(n608) );
  INV_X2 U2774 ( .A(n609), .ZN(n698) );
  INV_X2 U2775 ( .A(n602), .ZN(n600) );
  INV_X2 U2776 ( .A(n601), .ZN(n696) );
  INV_X2 U2777 ( .A(n594), .ZN(n592) );
  INV_X2 U2778 ( .A(n593), .ZN(n694) );
  INV_X2 U2779 ( .A(n586), .ZN(n584) );
  INV_X2 U2780 ( .A(n585), .ZN(n692) );
  INV_X2 U2781 ( .A(n578), .ZN(n576) );
  INV_X2 U2782 ( .A(n577), .ZN(n690) );
  INV_X2 U2783 ( .A(n570), .ZN(n568) );
  INV_X2 U2784 ( .A(n569), .ZN(n688) );
  INV_X2 U2785 ( .A(n562), .ZN(n560) );
  INV_X2 U2786 ( .A(n561), .ZN(n686) );
  INV_X2 U2787 ( .A(n554), .ZN(n552) );
  INV_X2 U2788 ( .A(n553), .ZN(n684) );
  INV_X2 U2789 ( .A(n390), .ZN(n2841) );
  INV_X2 U2790 ( .A(n2873), .ZN(n2839) );
  INV_X2 U2791 ( .A(n2872), .ZN(n2838) );
  INV_X2 U2792 ( .A(n2871), .ZN(n2837) );
  INV_X2 U2793 ( .A(n2870), .ZN(n2836) );
  INV_X2 U2794 ( .A(n2869), .ZN(n2835) );
  INV_X2 U2795 ( .A(n2868), .ZN(n2834) );
  INV_X2 U2796 ( .A(n2867), .ZN(n2833) );
  INV_X2 U2797 ( .A(n2866), .ZN(n2832) );
  INV_X2 U2798 ( .A(n2865), .ZN(n2831) );
  INV_X2 U2799 ( .A(n2864), .ZN(n2830) );
  INV_X2 U2800 ( .A(n2863), .ZN(n2829) );
  INV_X2 U2801 ( .A(n2862), .ZN(n2828) );
  INV_X2 U2802 ( .A(n2861), .ZN(n2827) );
  INV_X2 U2803 ( .A(n2860), .ZN(n2826) );
  INV_X2 U2804 ( .A(n2859), .ZN(n2825) );
  INV_X2 U2805 ( .A(n2858), .ZN(n2824) );
  INV_X2 U2806 ( .A(n2857), .ZN(n2823) );
  INV_X2 U2807 ( .A(n2856), .ZN(n2822) );
  INV_X2 U2808 ( .A(n2855), .ZN(n2821) );
  INV_X2 U2809 ( .A(n2854), .ZN(n2820) );
  INV_X2 U2810 ( .A(n2853), .ZN(n2819) );
  INV_X2 U2811 ( .A(n2852), .ZN(n2818) );
  INV_X2 U2812 ( .A(n2851), .ZN(n2817) );
  INV_X2 U2813 ( .A(n2850), .ZN(n2816) );
  INV_X2 U2814 ( .A(n2849), .ZN(n2815) );
  INV_X2 U2815 ( .A(n2848), .ZN(n2814) );
  INV_X2 U2816 ( .A(n2847), .ZN(n2813) );
  INV_X2 U2817 ( .A(n2846), .ZN(n2812) );
  INV_X2 U2818 ( .A(n2845), .ZN(n2811) );
  INV_X2 U2819 ( .A(n2844), .ZN(n2810) );
  INV_X2 U2820 ( .A(n2843), .ZN(n2809) );
  INV_X2 U2821 ( .A(n1406), .ZN(n2807) );
  AOI22_X2 U2822 ( .A1(n3154), .A2(n393), .B1(n313), .B2(n390), .ZN(n2806) );
  INV_X2 U2823 ( .A(n3238), .ZN(n313) );
  INV_X2 U2824 ( .A(n1403), .ZN(n2739) );
  OR2_X2 U2825 ( .A1(n2928), .A2(n3237), .ZN(n3239) );
  INV_X2 U2826 ( .A(n2917), .ZN(n3237) );
  INV_X2 U2827 ( .A(n1400), .ZN(n2671) );
  AOI22_X2 U2828 ( .A1(n295), .A2(n393), .B1(n317), .B2(n390), .ZN(n2670) );
  OR2_X2 U2829 ( .A1(n2927), .A2(n3236), .ZN(n3240) );
  INV_X2 U2830 ( .A(n2916), .ZN(n3236) );
  INV_X2 U2831 ( .A(n1397), .ZN(n2603) );
  AOI22_X2 U2832 ( .A1(n297), .A2(n393), .B1(n319), .B2(n390), .ZN(n2602) );
  INV_X2 U2833 ( .A(n2915), .ZN(n3235) );
  INV_X2 U2834 ( .A(n1394), .ZN(n2535) );
  AOI22_X2 U2835 ( .A1(n3185), .A2(n393), .B1(n321), .B2(n390), .ZN(n2534) );
  INV_X2 U2836 ( .A(n3242), .ZN(n321) );
  OR2_X2 U2837 ( .A1(n2925), .A2(n3234), .ZN(n3242) );
  INV_X2 U2838 ( .A(n1391), .ZN(n2467) );
  AOI22_X2 U2839 ( .A1(n3142), .A2(n393), .B1(n323), .B2(n390), .ZN(n2466) );
  INV_X2 U2840 ( .A(n3243), .ZN(n323) );
  OR2_X2 U2841 ( .A1(n2924), .A2(n3233), .ZN(n3243) );
  INV_X2 U2842 ( .A(n2913), .ZN(n3233) );
  INV_X2 U2843 ( .A(n1388), .ZN(n2399) );
  AOI22_X2 U2844 ( .A1(n3139), .A2(n393), .B1(n325), .B2(n390), .ZN(n2398) );
  INV_X2 U2845 ( .A(n3244), .ZN(n325) );
  OR2_X2 U2846 ( .A1(n2923), .A2(n3232), .ZN(n3244) );
  INV_X2 U2847 ( .A(n2912), .ZN(n3232) );
  INV_X2 U2848 ( .A(n1385), .ZN(n2331) );
  AOI22_X2 U2849 ( .A1(n3136), .A2(n393), .B1(n327), .B2(n390), .ZN(n2330) );
  INV_X2 U2850 ( .A(n3245), .ZN(n327) );
  OR2_X2 U2851 ( .A1(n2922), .A2(n3231), .ZN(n3245) );
  INV_X2 U2852 ( .A(n2911), .ZN(n3231) );
  INV_X2 U2853 ( .A(n1382), .ZN(n2263) );
  AOI22_X2 U2854 ( .A1(n3151), .A2(n393), .B1(n329), .B2(n390), .ZN(n2262) );
  INV_X2 U2855 ( .A(n3246), .ZN(n329) );
  OR2_X2 U2856 ( .A1(n2921), .A2(n3230), .ZN(n3246) );
  INV_X2 U2857 ( .A(n2910), .ZN(n3230) );
  INV_X2 U2858 ( .A(n1379), .ZN(n2195) );
  AOI22_X2 U2859 ( .A1(n3148), .A2(n393), .B1(n331), .B2(n390), .ZN(n2194) );
  INV_X2 U2860 ( .A(n3247), .ZN(n331) );
  OR2_X2 U2861 ( .A1(n2920), .A2(n3229), .ZN(n3247) );
  INV_X2 U2862 ( .A(n2909), .ZN(n3229) );
  INV_X2 U2863 ( .A(n1376), .ZN(n2127) );
  AOI22_X2 U2864 ( .A1(n3144), .A2(n393), .B1(n333), .B2(n390), .ZN(n2126) );
  INV_X2 U2865 ( .A(n3248), .ZN(n333) );
  OR2_X2 U2866 ( .A1(n2919), .A2(n3228), .ZN(n3248) );
  INV_X2 U2867 ( .A(n2908), .ZN(n3228) );
  INV_X2 U2868 ( .A(n262), .ZN(n2059) );
  INV_X2 U2869 ( .A(n265), .ZN(n2024) );
  INV_X2 U2870 ( .A(n268), .ZN(n1989) );
  INV_X2 U2871 ( .A(n274), .ZN(n1919) );
  INV_X2 U2872 ( .A(n277), .ZN(n1884) );
  INV_X2 U2873 ( .A(n280), .ZN(n1849) );
  INV_X2 U2874 ( .A(n283), .ZN(n1814) );
  INV_X2 U2875 ( .A(n286), .ZN(n1779) );
  INV_X2 U2876 ( .A(n289), .ZN(n1745) );
  INV_X2 U2877 ( .A(n1686), .ZN(n1719) );
  INV_X2 U2878 ( .A(n1682), .ZN(n1718) );
  INV_X2 U2879 ( .A(n1679), .ZN(n1717) );
  INV_X2 U2880 ( .A(n1668), .ZN(n1715) );
  INV_X2 U2881 ( .A(n1663), .ZN(n1714) );
  INV_X2 U2882 ( .A(n1660), .ZN(n1713) );
  INV_X2 U2883 ( .A(n1652), .ZN(n1712) );
  INV_X2 U2884 ( .A(n1649), .ZN(n1711) );
  INV_X2 U2885 ( .A(n1637), .ZN(n1709) );
  INV_X2 U2886 ( .A(n1621), .ZN(n1707) );
  INV_X2 U2887 ( .A(n1607), .ZN(n1705) );
  INV_X2 U2888 ( .A(n1592), .ZN(n1703) );
  INV_X2 U2889 ( .A(n1581), .ZN(n1702) );
  INV_X2 U2890 ( .A(n1576), .ZN(n1701) );
  INV_X2 U2891 ( .A(n1561), .ZN(n1700) );
  INV_X2 U2892 ( .A(n1556), .ZN(n1699) );
  INV_X2 U2893 ( .A(n1543), .ZN(n1698) );
  INV_X2 U2894 ( .A(n1538), .ZN(n1697) );
  INV_X2 U2895 ( .A(n1523), .ZN(n1696) );
  INV_X2 U2896 ( .A(n1518), .ZN(n1695) );
  INV_X2 U2897 ( .A(n1496), .ZN(n1693) );
  INV_X2 U2898 ( .A(n1474), .ZN(n1691) );
  INV_X2 U2899 ( .A(n1459), .ZN(n1690) );
  INV_X2 U2900 ( .A(n1450), .ZN(n1689) );
  INV_X2 U2901 ( .A(n1684), .ZN(n1685) );
  INV_X2 U2902 ( .A(n1676), .ZN(n1675) );
  INV_X2 U2903 ( .A(n1674), .ZN(n1672) );
  INV_X2 U2904 ( .A(n1673), .ZN(n1716) );
  INV_X2 U2905 ( .A(n1655), .ZN(n1654) );
  INV_X2 U2906 ( .A(n1648), .ZN(n1646) );
  INV_X2 U2907 ( .A(n1647), .ZN(n1645) );
  INV_X2 U2908 ( .A(n1643), .ZN(n1641) );
  INV_X2 U2909 ( .A(n1642), .ZN(n1710) );
  INV_X2 U2910 ( .A(n1630), .ZN(n1632) );
  INV_X2 U2911 ( .A(n1629), .ZN(n1631) );
  INV_X2 U2912 ( .A(n1627), .ZN(n1625) );
  INV_X2 U2913 ( .A(n1626), .ZN(n1708) );
  INV_X2 U2914 ( .A(n1613), .ZN(n1611) );
  INV_X2 U2915 ( .A(n1612), .ZN(n1706) );
  INV_X2 U2916 ( .A(n1600), .ZN(n1599) );
  INV_X2 U2917 ( .A(n1598), .ZN(n1596) );
  INV_X2 U2918 ( .A(n1597), .ZN(n1704) );
  INV_X2 U2919 ( .A(n1587), .ZN(n1589) );
  INV_X2 U2920 ( .A(n1586), .ZN(n1588) );
  INV_X2 U2921 ( .A(n1569), .ZN(n1571) );
  INV_X2 U2922 ( .A(n1568), .ZN(n1570) );
  INV_X2 U2923 ( .A(n1551), .ZN(n1549) );
  INV_X2 U2924 ( .A(n1550), .ZN(n1548) );
  INV_X2 U2925 ( .A(n1529), .ZN(n1531) );
  INV_X2 U2926 ( .A(n1528), .ZN(n1530) );
  INV_X2 U2927 ( .A(n1513), .ZN(n1511) );
  INV_X2 U2928 ( .A(n1512), .ZN(n1510) );
  INV_X2 U2929 ( .A(n1506), .ZN(n1504) );
  INV_X2 U2930 ( .A(n1505), .ZN(n1694) );
  INV_X2 U2931 ( .A(n1489), .ZN(n1491) );
  INV_X2 U2932 ( .A(n1488), .ZN(n1490) );
  INV_X2 U2933 ( .A(n1484), .ZN(n1482) );
  INV_X2 U2934 ( .A(n1483), .ZN(n1692) );
  INV_X2 U2935 ( .A(n1469), .ZN(n1471) );
  INV_X2 U2936 ( .A(n1468), .ZN(n1470) );
  INV_X2 U2937 ( .A(n484), .ZN(n1440) );
endmodule


module reg64_2 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  DFFR_X1 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module reg64_1 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  DFFR_X1 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module reg64_0 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  DFFR_X1 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module mul32_2 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_2_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module mul32_1 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_1_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module mul32_0 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_0_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module reg64_3 ( d, resetn, clk, q );
  input [63:0] d;
  output [63:0] q;
  input resetn, clk;
  wire   n65, n66, n67, n68, n69, n70;

  DFFR_X1 \q_reg[63]  ( .D(d[63]), .CK(clk), .RN(n70), .Q(q[63]) );
  DFFR_X1 \q_reg[62]  ( .D(d[62]), .CK(clk), .RN(n70), .Q(q[62]) );
  DFFR_X1 \q_reg[61]  ( .D(d[61]), .CK(clk), .RN(n70), .Q(q[61]) );
  DFFR_X1 \q_reg[60]  ( .D(d[60]), .CK(clk), .RN(n70), .Q(q[60]) );
  DFFR_X1 \q_reg[59]  ( .D(d[59]), .CK(clk), .RN(n69), .Q(q[59]) );
  DFFR_X1 \q_reg[58]  ( .D(d[58]), .CK(clk), .RN(n69), .Q(q[58]) );
  DFFR_X1 \q_reg[57]  ( .D(d[57]), .CK(clk), .RN(n69), .Q(q[57]) );
  DFFR_X1 \q_reg[56]  ( .D(d[56]), .CK(clk), .RN(n69), .Q(q[56]) );
  DFFR_X1 \q_reg[55]  ( .D(d[55]), .CK(clk), .RN(n69), .Q(q[55]) );
  DFFR_X1 \q_reg[54]  ( .D(d[54]), .CK(clk), .RN(n69), .Q(q[54]) );
  DFFR_X1 \q_reg[53]  ( .D(d[53]), .CK(clk), .RN(n69), .Q(q[53]) );
  DFFR_X1 \q_reg[52]  ( .D(d[52]), .CK(clk), .RN(n69), .Q(q[52]) );
  DFFR_X1 \q_reg[51]  ( .D(d[51]), .CK(clk), .RN(n69), .Q(q[51]) );
  DFFR_X1 \q_reg[50]  ( .D(d[50]), .CK(clk), .RN(n69), .Q(q[50]) );
  DFFR_X1 \q_reg[49]  ( .D(d[49]), .CK(clk), .RN(n69), .Q(q[49]) );
  DFFR_X1 \q_reg[48]  ( .D(d[48]), .CK(clk), .RN(n69), .Q(q[48]) );
  DFFR_X1 \q_reg[47]  ( .D(d[47]), .CK(clk), .RN(n68), .Q(q[47]) );
  DFFR_X1 \q_reg[46]  ( .D(d[46]), .CK(clk), .RN(n68), .Q(q[46]) );
  DFFR_X1 \q_reg[45]  ( .D(d[45]), .CK(clk), .RN(n68), .Q(q[45]) );
  DFFR_X1 \q_reg[44]  ( .D(d[44]), .CK(clk), .RN(n68), .Q(q[44]) );
  DFFR_X1 \q_reg[43]  ( .D(d[43]), .CK(clk), .RN(n68), .Q(q[43]) );
  DFFR_X1 \q_reg[42]  ( .D(d[42]), .CK(clk), .RN(n68), .Q(q[42]) );
  DFFR_X1 \q_reg[41]  ( .D(d[41]), .CK(clk), .RN(n68), .Q(q[41]) );
  DFFR_X1 \q_reg[40]  ( .D(d[40]), .CK(clk), .RN(n68), .Q(q[40]) );
  DFFR_X1 \q_reg[39]  ( .D(d[39]), .CK(clk), .RN(n68), .Q(q[39]) );
  DFFR_X1 \q_reg[38]  ( .D(d[38]), .CK(clk), .RN(n68), .Q(q[38]) );
  DFFR_X1 \q_reg[37]  ( .D(d[37]), .CK(clk), .RN(n68), .Q(q[37]) );
  DFFR_X1 \q_reg[36]  ( .D(d[36]), .CK(clk), .RN(n68), .Q(q[36]) );
  DFFR_X1 \q_reg[35]  ( .D(d[35]), .CK(clk), .RN(n67), .Q(q[35]) );
  DFFR_X1 \q_reg[34]  ( .D(d[34]), .CK(clk), .RN(n67), .Q(q[34]) );
  DFFR_X1 \q_reg[33]  ( .D(d[33]), .CK(clk), .RN(n67), .Q(q[33]) );
  DFFR_X1 \q_reg[32]  ( .D(d[32]), .CK(clk), .RN(n67), .Q(q[32]) );
  DFFR_X1 \q_reg[31]  ( .D(d[31]), .CK(clk), .RN(n67), .Q(q[31]) );
  DFFR_X1 \q_reg[30]  ( .D(d[30]), .CK(clk), .RN(n67), .Q(q[30]) );
  DFFR_X1 \q_reg[29]  ( .D(d[29]), .CK(clk), .RN(n67), .Q(q[29]) );
  DFFR_X1 \q_reg[28]  ( .D(d[28]), .CK(clk), .RN(n67), .Q(q[28]) );
  DFFR_X1 \q_reg[27]  ( .D(d[27]), .CK(clk), .RN(n67), .Q(q[27]) );
  DFFR_X1 \q_reg[26]  ( .D(d[26]), .CK(clk), .RN(n67), .Q(q[26]) );
  DFFR_X1 \q_reg[25]  ( .D(d[25]), .CK(clk), .RN(n67), .Q(q[25]) );
  DFFR_X1 \q_reg[24]  ( .D(d[24]), .CK(clk), .RN(n67), .Q(q[24]) );
  DFFR_X1 \q_reg[23]  ( .D(d[23]), .CK(clk), .RN(n66), .Q(q[23]) );
  DFFR_X1 \q_reg[22]  ( .D(d[22]), .CK(clk), .RN(n66), .Q(q[22]) );
  DFFR_X1 \q_reg[21]  ( .D(d[21]), .CK(clk), .RN(n66), .Q(q[21]) );
  DFFR_X1 \q_reg[20]  ( .D(d[20]), .CK(clk), .RN(n66), .Q(q[20]) );
  DFFR_X1 \q_reg[19]  ( .D(d[19]), .CK(clk), .RN(n66), .Q(q[19]) );
  DFFR_X1 \q_reg[18]  ( .D(d[18]), .CK(clk), .RN(n66), .Q(q[18]) );
  DFFR_X1 \q_reg[17]  ( .D(d[17]), .CK(clk), .RN(n66), .Q(q[17]) );
  DFFR_X1 \q_reg[16]  ( .D(d[16]), .CK(clk), .RN(n66), .Q(q[16]) );
  DFFR_X1 \q_reg[15]  ( .D(d[15]), .CK(clk), .RN(n66), .Q(q[15]) );
  DFFR_X1 \q_reg[14]  ( .D(d[14]), .CK(clk), .RN(n66), .Q(q[14]) );
  DFFR_X1 \q_reg[13]  ( .D(d[13]), .CK(clk), .RN(n66), .Q(q[13]) );
  DFFR_X1 \q_reg[12]  ( .D(d[12]), .CK(clk), .RN(n66), .Q(q[12]) );
  DFFR_X1 \q_reg[11]  ( .D(d[11]), .CK(clk), .RN(n65), .Q(q[11]) );
  DFFR_X1 \q_reg[10]  ( .D(d[10]), .CK(clk), .RN(n65), .Q(q[10]) );
  DFFR_X1 \q_reg[9]  ( .D(d[9]), .CK(clk), .RN(n65), .Q(q[9]) );
  DFFR_X1 \q_reg[8]  ( .D(d[8]), .CK(clk), .RN(n65), .Q(q[8]) );
  DFFR_X1 \q_reg[7]  ( .D(d[7]), .CK(clk), .RN(n65), .Q(q[7]) );
  DFFR_X1 \q_reg[6]  ( .D(d[6]), .CK(clk), .RN(n65), .Q(q[6]) );
  DFFR_X1 \q_reg[5]  ( .D(d[5]), .CK(clk), .RN(n65), .Q(q[5]) );
  DFFR_X1 \q_reg[4]  ( .D(d[4]), .CK(clk), .RN(n65), .Q(q[4]) );
  DFFR_X1 \q_reg[3]  ( .D(d[3]), .CK(clk), .RN(n65), .Q(q[3]) );
  DFFR_X1 \q_reg[2]  ( .D(d[2]), .CK(clk), .RN(n65), .Q(q[2]) );
  DFFR_X1 \q_reg[1]  ( .D(d[1]), .CK(clk), .RN(n65), .Q(q[1]) );
  DFFR_X1 \q_reg[0]  ( .D(d[0]), .CK(clk), .RN(n65), .Q(q[0]) );
  BUF_X1 U3 ( .A(resetn), .Z(n65) );
  BUF_X1 U4 ( .A(resetn), .Z(n66) );
  BUF_X1 U5 ( .A(resetn), .Z(n67) );
  BUF_X1 U6 ( .A(resetn), .Z(n68) );
  BUF_X1 U7 ( .A(resetn), .Z(n69) );
  BUF_X1 U8 ( .A(resetn), .Z(n70) );
endmodule


module mul32_3 ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;


  mul32_3_DW_mult_uns_1 mult_12 ( .a(a), .b(b), .product(result) );
endmodule


module mulcascade ( a0, b0, a1, b1, a2, b2, a3, b3, result0, result1, result2, 
        result3, resetn, clk );
  input [31:0] a0;
  input [31:0] b0;
  input [31:0] a1;
  input [31:0] b1;
  input [31:0] a2;
  input [31:0] b2;
  input [31:0] a3;
  input [31:0] b3;
  output [63:0] result0;
  output [63:0] result1;
  output [63:0] result2;
  output [63:0] result3;
  input resetn, clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173;
  wire   [63:0] reg0in;
  wire   [63:0] reg1in;
  wire   [63:0] reg2in;
  wire   [63:0] reg3in;

  mul32_3 mul0 ( .a({n89, n27, n170, n11, n22, n171, n23, n34, n172, n39, n26, 
        a0[20], n30, n18, a0[17], n19, n76, a0[14], n81, n52, a0[11], n69, n60, 
        a0[8], n47, n42, a0[5], n38, n35, a0[2], n31, n88}), .b({n130, n128, 
        n129, n133, n126, n127, n158, n161, n155, n156, n150, n153, n147, n148, 
        n142, n145, b0[15:1], n91}), .result(reg0in) );
  reg64_3 reg0 ( .d(reg0in), .resetn(n173), .clk(clk), .q(result0) );
  mul32_2 mul1 ( .a({n85, n15, n165, n14, n10, n166, n7, n6, a1[23], n3, n2, 
        a1[20], n80, n77, a1[17], n73, n72, a1[14], n68, n65, a1[11], n64, n61, 
        a1[8], n57, n55, a1[5], n51, n48, a1[2], n44, n84}), .b({n124, n125, 
        n123, n122, n120, n121, n118, n117, n113, n116, n111, n110, n105, n108, 
        n103, n102, b1[15:0]}), .result(reg1in) );
  reg64_2 reg1 ( .d(reg1in), .resetn(n173), .clk(clk), .q(result1) );
  mul32_1 mul2 ( .a({n86, n4, n162, n8, n9, n164, n12, n13, n163, n17, n20, 
        a2[20], n21, n24, a2[17], n28, n29, a2[14], n33, n36, a2[11], n40, n41, 
        a2[8], n45, n46, a2[5], n50, n53, a2[2], n58, n87}), .b({n95, n94, n96, 
        n97, n99, n98, n100, n101, n106, n104, n107, n109, n114, n112, n115, 
        n119, b2[15:0]}), .result(reg2in) );
  reg64_1 reg2 ( .d(reg2in), .resetn(n173), .clk(clk), .q(result2) );
  mul32_0 mul3 ( .a({n83, n71, n167, n74, n78, n168, n79, n1, n169, n5, n25, 
        a3[20], n16, n37, a3[17], n32, n59, a3[14], n54, n66, a3[11], n63, n70, 
        a3[8], n82, n75, a3[5], n67, n62, a3[2], n49, n90}), .b({n136, n138, 
        n137, n139, n140, n141, n143, n144, n146, n149, n151, n152, n154, n157, 
        n159, n160, n135, n132, n93, n131, b3[11:0]}), .result(reg3in) );
  reg64_0 reg4 ( .d(reg3in), .resetn(n173), .clk(clk), .q(result3) );
  BUF_X4 U1 ( .A(b3[12]), .Z(n131) );
  BUF_X4 U2 ( .A(b3[14]), .Z(n132) );
  INV_X1 U3 ( .A(b3[15]), .ZN(n134) );
  INV_X1 U4 ( .A(b3[13]), .ZN(n92) );
  BUF_X1 U5 ( .A(a3[24]), .Z(n1) );
  BUF_X1 U6 ( .A(a1[21]), .Z(n2) );
  BUF_X1 U7 ( .A(a1[22]), .Z(n3) );
  BUF_X1 U8 ( .A(a2[30]), .Z(n4) );
  BUF_X1 U9 ( .A(a3[22]), .Z(n5) );
  BUF_X1 U10 ( .A(a1[24]), .Z(n6) );
  BUF_X1 U11 ( .A(a1[25]), .Z(n7) );
  BUF_X1 U12 ( .A(a2[28]), .Z(n8) );
  BUF_X1 U13 ( .A(a2[27]), .Z(n9) );
  BUF_X1 U14 ( .A(a1[27]), .Z(n10) );
  BUF_X1 U15 ( .A(a0[28]), .Z(n11) );
  BUF_X1 U16 ( .A(a2[25]), .Z(n12) );
  BUF_X1 U17 ( .A(a2[24]), .Z(n13) );
  BUF_X1 U18 ( .A(a1[28]), .Z(n14) );
  BUF_X1 U19 ( .A(a1[30]), .Z(n15) );
  BUF_X1 U20 ( .A(a3[19]), .Z(n16) );
  BUF_X1 U21 ( .A(a2[22]), .Z(n17) );
  BUF_X1 U22 ( .A(a0[18]), .Z(n18) );
  BUF_X1 U23 ( .A(a0[16]), .Z(n19) );
  BUF_X1 U24 ( .A(a2[21]), .Z(n20) );
  BUF_X1 U25 ( .A(a2[19]), .Z(n21) );
  BUF_X1 U26 ( .A(a0[27]), .Z(n22) );
  BUF_X1 U27 ( .A(a0[25]), .Z(n23) );
  BUF_X1 U28 ( .A(a2[18]), .Z(n24) );
  BUF_X1 U29 ( .A(a3[21]), .Z(n25) );
  BUF_X1 U30 ( .A(a0[21]), .Z(n26) );
  BUF_X1 U31 ( .A(a0[30]), .Z(n27) );
  BUF_X1 U32 ( .A(a2[16]), .Z(n28) );
  BUF_X1 U33 ( .A(a2[15]), .Z(n29) );
  BUF_X1 U34 ( .A(a0[19]), .Z(n30) );
  BUF_X1 U35 ( .A(a0[1]), .Z(n31) );
  BUF_X1 U36 ( .A(a3[16]), .Z(n32) );
  BUF_X1 U37 ( .A(a2[13]), .Z(n33) );
  BUF_X1 U38 ( .A(a0[24]), .Z(n34) );
  BUF_X1 U39 ( .A(a0[3]), .Z(n35) );
  BUF_X1 U40 ( .A(a2[12]), .Z(n36) );
  BUF_X1 U41 ( .A(a3[18]), .Z(n37) );
  BUF_X1 U42 ( .A(a0[4]), .Z(n38) );
  BUF_X1 U43 ( .A(a0[22]), .Z(n39) );
  BUF_X1 U44 ( .A(a2[10]), .Z(n40) );
  BUF_X1 U45 ( .A(a2[9]), .Z(n41) );
  BUF_X1 U46 ( .A(a0[6]), .Z(n42) );
  INV_X1 U47 ( .A(a1[1]), .ZN(n43) );
  INV_X1 U48 ( .A(n43), .ZN(n44) );
  BUF_X1 U49 ( .A(a2[7]), .Z(n45) );
  BUF_X1 U50 ( .A(a2[6]), .Z(n46) );
  BUF_X1 U51 ( .A(a0[7]), .Z(n47) );
  BUF_X1 U52 ( .A(a1[3]), .Z(n48) );
  BUF_X1 U53 ( .A(a3[1]), .Z(n49) );
  BUF_X1 U54 ( .A(a2[4]), .Z(n50) );
  BUF_X1 U55 ( .A(a1[4]), .Z(n51) );
  BUF_X1 U56 ( .A(a0[12]), .Z(n52) );
  BUF_X1 U57 ( .A(a2[3]), .Z(n53) );
  BUF_X1 U58 ( .A(a3[13]), .Z(n54) );
  BUF_X2 U59 ( .A(a1[6]), .Z(n55) );
  INV_X1 U60 ( .A(a1[7]), .ZN(n56) );
  INV_X1 U61 ( .A(n56), .ZN(n57) );
  BUF_X1 U62 ( .A(a2[1]), .Z(n58) );
  BUF_X1 U63 ( .A(a3[15]), .Z(n59) );
  BUF_X1 U64 ( .A(a0[9]), .Z(n60) );
  BUF_X1 U65 ( .A(a1[9]), .Z(n61) );
  BUF_X1 U66 ( .A(a3[3]), .Z(n62) );
  BUF_X1 U67 ( .A(a3[10]), .Z(n63) );
  BUF_X2 U68 ( .A(a1[10]), .Z(n64) );
  BUF_X1 U69 ( .A(a1[12]), .Z(n65) );
  BUF_X1 U70 ( .A(a3[12]), .Z(n66) );
  BUF_X1 U71 ( .A(a3[4]), .Z(n67) );
  BUF_X1 U72 ( .A(a1[13]), .Z(n68) );
  BUF_X1 U73 ( .A(a0[10]), .Z(n69) );
  BUF_X1 U74 ( .A(a3[9]), .Z(n70) );
  BUF_X1 U75 ( .A(a3[30]), .Z(n71) );
  BUF_X1 U76 ( .A(a1[15]), .Z(n72) );
  BUF_X1 U77 ( .A(a1[16]), .Z(n73) );
  BUF_X1 U78 ( .A(a3[28]), .Z(n74) );
  BUF_X1 U79 ( .A(a3[6]), .Z(n75) );
  BUF_X1 U80 ( .A(a0[15]), .Z(n76) );
  BUF_X1 U81 ( .A(a1[18]), .Z(n77) );
  BUF_X1 U82 ( .A(a3[27]), .Z(n78) );
  BUF_X1 U83 ( .A(a3[25]), .Z(n79) );
  BUF_X1 U84 ( .A(a1[19]), .Z(n80) );
  BUF_X1 U85 ( .A(a0[13]), .Z(n81) );
  BUF_X1 U86 ( .A(a3[7]), .Z(n82) );
  BUF_X1 U87 ( .A(a3[31]), .Z(n83) );
  BUF_X1 U88 ( .A(a1[0]), .Z(n84) );
  BUF_X1 U89 ( .A(a1[31]), .Z(n85) );
  BUF_X1 U90 ( .A(a2[31]), .Z(n86) );
  BUF_X1 U91 ( .A(a2[0]), .Z(n87) );
  BUF_X1 U92 ( .A(a0[0]), .Z(n88) );
  BUF_X1 U93 ( .A(a0[31]), .Z(n89) );
  BUF_X1 U94 ( .A(a3[0]), .Z(n90) );
  BUF_X4 U95 ( .A(b0[0]), .Z(n91) );
  INV_X4 U96 ( .A(n92), .ZN(n93) );
  BUF_X4 U97 ( .A(b2[30]), .Z(n94) );
  BUF_X4 U98 ( .A(b2[31]), .Z(n95) );
  BUF_X4 U99 ( .A(b2[29]), .Z(n96) );
  BUF_X4 U100 ( .A(b2[28]), .Z(n97) );
  BUF_X4 U101 ( .A(b2[26]), .Z(n98) );
  BUF_X4 U102 ( .A(b2[27]), .Z(n99) );
  BUF_X4 U103 ( .A(b2[25]), .Z(n100) );
  BUF_X4 U104 ( .A(b2[24]), .Z(n101) );
  BUF_X4 U105 ( .A(b1[16]), .Z(n102) );
  BUF_X4 U106 ( .A(b1[17]), .Z(n103) );
  BUF_X4 U107 ( .A(b2[22]), .Z(n104) );
  BUF_X4 U108 ( .A(b1[19]), .Z(n105) );
  BUF_X4 U109 ( .A(b2[23]), .Z(n106) );
  BUF_X4 U110 ( .A(b2[21]), .Z(n107) );
  BUF_X4 U111 ( .A(b1[18]), .Z(n108) );
  BUF_X4 U112 ( .A(b2[20]), .Z(n109) );
  BUF_X4 U113 ( .A(b1[20]), .Z(n110) );
  BUF_X4 U114 ( .A(b1[21]), .Z(n111) );
  BUF_X4 U115 ( .A(b2[18]), .Z(n112) );
  BUF_X4 U116 ( .A(b1[23]), .Z(n113) );
  BUF_X4 U117 ( .A(b2[19]), .Z(n114) );
  BUF_X4 U118 ( .A(b2[17]), .Z(n115) );
  BUF_X4 U119 ( .A(b1[22]), .Z(n116) );
  BUF_X4 U120 ( .A(b1[24]), .Z(n117) );
  BUF_X4 U121 ( .A(b1[25]), .Z(n118) );
  BUF_X4 U122 ( .A(b2[16]), .Z(n119) );
  BUF_X4 U123 ( .A(b1[27]), .Z(n120) );
  BUF_X4 U124 ( .A(b1[26]), .Z(n121) );
  BUF_X4 U125 ( .A(b1[28]), .Z(n122) );
  BUF_X4 U126 ( .A(b1[29]), .Z(n123) );
  BUF_X4 U127 ( .A(b1[31]), .Z(n124) );
  BUF_X4 U128 ( .A(b1[30]), .Z(n125) );
  BUF_X4 U129 ( .A(b0[27]), .Z(n126) );
  BUF_X4 U130 ( .A(b0[26]), .Z(n127) );
  BUF_X4 U131 ( .A(b0[30]), .Z(n128) );
  BUF_X4 U132 ( .A(b0[29]), .Z(n129) );
  BUF_X4 U133 ( .A(b0[31]), .Z(n130) );
  BUF_X4 U134 ( .A(b0[28]), .Z(n133) );
  INV_X4 U135 ( .A(n134), .ZN(n135) );
  BUF_X4 U136 ( .A(b3[31]), .Z(n136) );
  BUF_X4 U137 ( .A(b3[29]), .Z(n137) );
  BUF_X4 U138 ( .A(b3[30]), .Z(n138) );
  BUF_X4 U139 ( .A(b3[28]), .Z(n139) );
  BUF_X4 U140 ( .A(b3[27]), .Z(n140) );
  BUF_X4 U141 ( .A(b3[26]), .Z(n141) );
  BUF_X4 U142 ( .A(b0[17]), .Z(n142) );
  BUF_X4 U143 ( .A(b3[25]), .Z(n143) );
  BUF_X4 U144 ( .A(b3[24]), .Z(n144) );
  BUF_X4 U145 ( .A(b0[16]), .Z(n145) );
  BUF_X4 U146 ( .A(b3[23]), .Z(n146) );
  BUF_X4 U147 ( .A(b0[19]), .Z(n147) );
  BUF_X4 U148 ( .A(b0[18]), .Z(n148) );
  BUF_X4 U149 ( .A(b3[22]), .Z(n149) );
  BUF_X4 U150 ( .A(b0[21]), .Z(n150) );
  BUF_X4 U151 ( .A(b3[21]), .Z(n151) );
  BUF_X4 U152 ( .A(b3[20]), .Z(n152) );
  BUF_X4 U153 ( .A(b0[20]), .Z(n153) );
  BUF_X4 U154 ( .A(b3[19]), .Z(n154) );
  BUF_X4 U155 ( .A(b0[23]), .Z(n155) );
  BUF_X4 U156 ( .A(b0[22]), .Z(n156) );
  BUF_X4 U157 ( .A(b3[18]), .Z(n157) );
  BUF_X4 U158 ( .A(b0[25]), .Z(n158) );
  BUF_X4 U159 ( .A(b3[17]), .Z(n159) );
  BUF_X4 U160 ( .A(b3[16]), .Z(n160) );
  BUF_X4 U161 ( .A(b0[24]), .Z(n161) );
  BUF_X4 U162 ( .A(a2[29]), .Z(n162) );
  BUF_X4 U163 ( .A(a2[23]), .Z(n163) );
  BUF_X4 U164 ( .A(a2[26]), .Z(n164) );
  BUF_X4 U165 ( .A(a1[29]), .Z(n165) );
  BUF_X4 U166 ( .A(a1[26]), .Z(n166) );
  BUF_X4 U167 ( .A(a3[29]), .Z(n167) );
  BUF_X4 U168 ( .A(a3[26]), .Z(n168) );
  BUF_X4 U169 ( .A(a3[23]), .Z(n169) );
  BUF_X4 U170 ( .A(a0[29]), .Z(n170) );
  BUF_X4 U171 ( .A(a0[26]), .Z(n171) );
  BUF_X4 U172 ( .A(a0[23]), .Z(n172) );
  BUF_X2 U173 ( .A(resetn), .Z(n173) );
endmodule

